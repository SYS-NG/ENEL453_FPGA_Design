LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY buzzer IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;		                         
      distance       :  IN    STD_LOGIC_VECTOR(12 DOWNTO 0);
		dac_out        :  OUT   STD_LOGIC
		);
END buzzer;

ARCHITECTURE behavior OF buzzer IS

signal counter       : unsigned(17 DOWNTO 0) := (others=>'0');
signal counter_limit : unsigned(17 DOWNTO 0);

type array_1d is array (0 to 4095) of integer;
	
constant d2count: array_1d := (
(	16519	)	,
(	16527	)	,
(	16535	)	,
(	16543	)	,
(	16551	)	,
(	16559	)	,
(	16567	)	,
(	16575	)	,
(	16582	)	,
(	16590	)	,
(	16598	)	,
(	16606	)	,
(	16614	)	,
(	16622	)	,
(	16630	)	,
(	16638	)	,
(	16646	)	,
(	16654	)	,
(	16662	)	,
(	16670	)	,
(	16678	)	,
(	16686	)	,
(	16694	)	,
(	16702	)	,
(	16710	)	,
(	16718	)	,
(	16726	)	,
(	16734	)	,
(	16742	)	,
(	16750	)	,
(	16758	)	,
(	16766	)	,
(	16774	)	,
(	16782	)	,
(	16790	)	,
(	16798	)	,
(	16806	)	,
(	16814	)	,
(	16822	)	,
(	16830	)	,
(	16838	)	,
(	16846	)	,
(	16854	)	,
(	16862	)	,
(	16870	)	,
(	16878	)	,
(	16886	)	,
(	16894	)	,
(	16903	)	,
(	16911	)	,
(	16919	)	,
(	16927	)	,
(	16935	)	,
(	16943	)	,
(	16951	)	,
(	16959	)	,
(	16967	)	,
(	16975	)	,
(	16984	)	,
(	16992	)	,
(	17000	)	,
(	17008	)	,
(	17016	)	,
(	17024	)	,
(	17032	)	,
(	17040	)	,
(	17049	)	,
(	17057	)	,
(	17065	)	,
(	17073	)	,
(	17081	)	,
(	17089	)	,
(	17098	)	,
(	17106	)	,
(	17114	)	,
(	17122	)	,
(	17130	)	,
(	17139	)	,
(	17147	)	,
(	17155	)	,
(	17163	)	,
(	17171	)	,
(	17180	)	,
(	17188	)	,
(	17196	)	,
(	17204	)	,
(	17212	)	,
(	17221	)	,
(	17229	)	,
(	17237	)	,
(	17245	)	,
(	17254	)	,
(	17262	)	,
(	17270	)	,
(	17278	)	,
(	17287	)	,
(	17295	)	,
(	17303	)	,
(	17311	)	,
(	17320	)	,
(	17328	)	,
(	17336	)	,
(	17345	)	,
(	17353	)	,
(	17361	)	,
(	17369	)	,
(	17378	)	,
(	17386	)	,
(	17394	)	,
(	17403	)	,
(	17411	)	,
(	17419	)	,
(	17428	)	,
(	17436	)	,
(	17444	)	,
(	17453	)	,
(	17461	)	,
(	17469	)	,
(	17478	)	,
(	17486	)	,
(	17494	)	,
(	17503	)	,
(	17511	)	,
(	17520	)	,
(	17528	)	,
(	17536	)	,
(	17545	)	,
(	17553	)	,
(	17561	)	,
(	17570	)	,
(	17578	)	,
(	17587	)	,
(	17595	)	,
(	17603	)	,
(	17612	)	,
(	17620	)	,
(	17629	)	,
(	17637	)	,
(	17646	)	,
(	17654	)	,
(	17663	)	,
(	17671	)	,
(	17679	)	,
(	17688	)	,
(	17696	)	,
(	17705	)	,
(	17713	)	,
(	17722	)	,
(	17730	)	,
(	17739	)	,
(	17747	)	,
(	17756	)	,
(	17764	)	,
(	17773	)	,
(	17781	)	,
(	17790	)	,
(	17798	)	,
(	17807	)	,
(	17815	)	,
(	17824	)	,
(	17832	)	,
(	17841	)	,
(	17849	)	,
(	17858	)	,
(	17866	)	,
(	17875	)	,
(	17883	)	,
(	17892	)	,
(	17901	)	,
(	17909	)	,
(	17918	)	,
(	17926	)	,
(	17935	)	,
(	17943	)	,
(	17952	)	,
(	17961	)	,
(	17969	)	,
(	17978	)	,
(	17986	)	,
(	17995	)	,
(	18003	)	,
(	18012	)	,
(	18021	)	,
(	18029	)	,
(	18038	)	,
(	18047	)	,
(	18055	)	,
(	18064	)	,
(	18072	)	,
(	18081	)	,
(	18090	)	,
(	18098	)	,
(	18107	)	,
(	18116	)	,
(	18124	)	,
(	18133	)	,
(	18142	)	,
(	18150	)	,
(	18159	)	,
(	18168	)	,
(	18176	)	,
(	18185	)	,
(	18194	)	,
(	18203	)	,
(	18211	)	,
(	18220	)	,
(	18229	)	,
(	18237	)	,
(	18246	)	,
(	18255	)	,
(	18264	)	,
(	18272	)	,
(	18281	)	,
(	18290	)	,
(	18298	)	,
(	18307	)	,
(	18316	)	,
(	18325	)	,
(	18334	)	,
(	18342	)	,
(	18351	)	,
(	18360	)	,
(	18369	)	,
(	18377	)	,
(	18386	)	,
(	18395	)	,
(	18404	)	,
(	18413	)	,
(	18421	)	,
(	18430	)	,
(	18439	)	,
(	18448	)	,
(	18457	)	,
(	18465	)	,
(	18474	)	,
(	18483	)	,
(	18492	)	,
(	18501	)	,
(	18510	)	,
(	18518	)	,
(	18527	)	,
(	18536	)	,
(	18545	)	,
(	18554	)	,
(	18563	)	,
(	18572	)	,
(	18581	)	,
(	18589	)	,
(	18598	)	,
(	18607	)	,
(	18616	)	,
(	18625	)	,
(	18634	)	,
(	18643	)	,
(	18652	)	,
(	18661	)	,
(	18670	)	,
(	18679	)	,
(	18687	)	,
(	18696	)	,
(	18705	)	,
(	18714	)	,
(	18723	)	,
(	18732	)	,
(	18741	)	,
(	18750	)	,
(	18759	)	,
(	18768	)	,
(	18777	)	,
(	18786	)	,
(	18795	)	,
(	18804	)	,
(	18813	)	,
(	18822	)	,
(	18831	)	,
(	18840	)	,
(	18849	)	,
(	18858	)	,
(	18867	)	,
(	18876	)	,
(	18885	)	,
(	18894	)	,
(	18903	)	,
(	18912	)	,
(	18921	)	,
(	18930	)	,
(	18939	)	,
(	18948	)	,
(	18957	)	,
(	18966	)	,
(	18976	)	,
(	18985	)	,
(	18994	)	,
(	19003	)	,
(	19012	)	,
(	19021	)	,
(	19030	)	,
(	19039	)	,
(	19048	)	,
(	19057	)	,
(	19066	)	,
(	19076	)	,
(	19085	)	,
(	19094	)	,
(	19103	)	,
(	19112	)	,
(	19121	)	,
(	19130	)	,
(	19139	)	,
(	19149	)	,
(	19158	)	,
(	19167	)	,
(	19176	)	,
(	19185	)	,
(	19194	)	,
(	19204	)	,
(	19213	)	,
(	19222	)	,
(	19231	)	,
(	19240	)	,
(	19250	)	,
(	19259	)	,
(	19268	)	,
(	19277	)	,
(	19286	)	,
(	19296	)	,
(	19305	)	,
(	19314	)	,
(	19323	)	,
(	19333	)	,
(	19342	)	,
(	19351	)	,
(	19360	)	,
(	19370	)	,
(	19379	)	,
(	19388	)	,
(	19397	)	,
(	19407	)	,
(	19416	)	,
(	19425	)	,
(	19435	)	,
(	19444	)	,
(	19453	)	,
(	19462	)	,
(	19472	)	,
(	19481	)	,
(	19490	)	,
(	19500	)	,
(	19509	)	,
(	19518	)	,
(	19528	)	,
(	19537	)	,
(	19546	)	,
(	19556	)	,
(	19565	)	,
(	19574	)	,
(	19584	)	,
(	19593	)	,
(	19602	)	,
(	19612	)	,
(	19621	)	,
(	19631	)	,
(	19640	)	,
(	19649	)	,
(	19659	)	,
(	19668	)	,
(	19678	)	,
(	19687	)	,
(	19696	)	,
(	19706	)	,
(	19715	)	,
(	19725	)	,
(	19734	)	,
(	19744	)	,
(	19753	)	,
(	19762	)	,
(	19772	)	,
(	19781	)	,
(	19791	)	,
(	19800	)	,
(	19810	)	,
(	19819	)	,
(	19829	)	,
(	19838	)	,
(	19848	)	,
(	19857	)	,
(	19867	)	,
(	19876	)	,
(	19886	)	,
(	19895	)	,
(	19905	)	,
(	19914	)	,
(	19924	)	,
(	19933	)	,
(	19943	)	,
(	19952	)	,
(	19962	)	,
(	19971	)	,
(	19981	)	,
(	19990	)	,
(	20000	)	,
(	20010	)	,
(	20019	)	,
(	20029	)	,
(	20038	)	,
(	20048	)	,
(	20057	)	,
(	20067	)	,
(	20077	)	,
(	20086	)	,
(	20096	)	,
(	20105	)	,
(	20115	)	,
(	20125	)	,
(	20134	)	,
(	20144	)	,
(	20154	)	,
(	20163	)	,
(	20173	)	,
(	20182	)	,
(	20192	)	,
(	20202	)	,
(	20211	)	,
(	20221	)	,
(	20231	)	,
(	20240	)	,
(	20250	)	,
(	20260	)	,
(	20269	)	,
(	20279	)	,
(	20289	)	,
(	20299	)	,
(	20308	)	,
(	20318	)	,
(	20328	)	,
(	20337	)	,
(	20347	)	,
(	20357	)	,
(	20367	)	,
(	20376	)	,
(	20386	)	,
(	20396	)	,
(	20406	)	,
(	20415	)	,
(	20425	)	,
(	20435	)	,
(	20445	)	,
(	20454	)	,
(	20464	)	,
(	20474	)	,
(	20484	)	,
(	20494	)	,
(	20503	)	,
(	20513	)	,
(	20523	)	,
(	20533	)	,
(	20543	)	,
(	20552	)	,
(	20562	)	,
(	20572	)	,
(	20582	)	,
(	20592	)	,
(	20602	)	,
(	20611	)	,
(	20621	)	,
(	20631	)	,
(	20641	)	,
(	20651	)	,
(	20661	)	,
(	20671	)	,
(	20681	)	,
(	20690	)	,
(	20700	)	,
(	20710	)	,
(	20720	)	,
(	20730	)	,
(	20740	)	,
(	20750	)	,
(	20760	)	,
(	20770	)	,
(	20780	)	,
(	20790	)	,
(	20800	)	,
(	20809	)	,
(	20819	)	,
(	20829	)	,
(	20839	)	,
(	20849	)	,
(	20859	)	,
(	20869	)	,
(	20879	)	,
(	20889	)	,
(	20899	)	,
(	20909	)	,
(	20919	)	,
(	20929	)	,
(	20939	)	,
(	20949	)	,
(	20959	)	,
(	20969	)	,
(	20979	)	,
(	20989	)	,
(	20999	)	,
(	21009	)	,
(	21019	)	,
(	21029	)	,
(	21040	)	,
(	21050	)	,
(	21060	)	,
(	21070	)	,
(	21080	)	,
(	21090	)	,
(	21100	)	,
(	21110	)	,
(	21120	)	,
(	21130	)	,
(	21140	)	,
(	21150	)	,
(	21161	)	,
(	21171	)	,
(	21181	)	,
(	21191	)	,
(	21201	)	,
(	21211	)	,
(	21221	)	,
(	21232	)	,
(	21242	)	,
(	21252	)	,
(	21262	)	,
(	21272	)	,
(	21282	)	,
(	21292	)	,
(	21303	)	,
(	21313	)	,
(	21323	)	,
(	21333	)	,
(	21343	)	,
(	21354	)	,
(	21364	)	,
(	21374	)	,
(	21384	)	,
(	21395	)	,
(	21405	)	,
(	21415	)	,
(	21425	)	,
(	21435	)	,
(	21446	)	,
(	21456	)	,
(	21466	)	,
(	21476	)	,
(	21487	)	,
(	21497	)	,
(	21507	)	,
(	21518	)	,
(	21528	)	,
(	21538	)	,
(	21548	)	,
(	21559	)	,
(	21569	)	,
(	21579	)	,
(	21590	)	,
(	21600	)	,
(	21610	)	,
(	21621	)	,
(	21631	)	,
(	21641	)	,
(	21652	)	,
(	21662	)	,
(	21672	)	,
(	21683	)	,
(	21693	)	,
(	21704	)	,
(	21714	)	,
(	21724	)	,
(	21735	)	,
(	21745	)	,
(	21755	)	,
(	21766	)	,
(	21776	)	,
(	21787	)	,
(	21797	)	,
(	21808	)	,
(	21818	)	,
(	21828	)	,
(	21839	)	,
(	21849	)	,
(	21860	)	,
(	21870	)	,
(	21881	)	,
(	21891	)	,
(	21902	)	,
(	21912	)	,
(	21923	)	,
(	21933	)	,
(	21943	)	,
(	21954	)	,
(	21964	)	,
(	21975	)	,
(	21985	)	,
(	21996	)	,
(	22007	)	,
(	22017	)	,
(	22028	)	,
(	22038	)	,
(	22049	)	,
(	22059	)	,
(	22070	)	,
(	22080	)	,
(	22091	)	,
(	22101	)	,
(	22112	)	,
(	22123	)	,
(	22133	)	,
(	22144	)	,
(	22154	)	,
(	22165	)	,
(	22175	)	,
(	22186	)	,
(	22197	)	,
(	22207	)	,
(	22218	)	,
(	22229	)	,
(	22239	)	,
(	22250	)	,
(	22260	)	,
(	22271	)	,
(	22282	)	,
(	22292	)	,
(	22303	)	,
(	22314	)	,
(	22324	)	,
(	22335	)	,
(	22346	)	,
(	22356	)	,
(	22367	)	,
(	22378	)	,
(	22389	)	,
(	22399	)	,
(	22410	)	,
(	22421	)	,
(	22431	)	,
(	22442	)	,
(	22453	)	,
(	22464	)	,
(	22474	)	,
(	22485	)	,
(	22496	)	,
(	22507	)	,
(	22517	)	,
(	22528	)	,
(	22539	)	,
(	22550	)	,
(	22560	)	,
(	22571	)	,
(	22582	)	,
(	22593	)	,
(	22604	)	,
(	22614	)	,
(	22625	)	,
(	22636	)	,
(	22647	)	,
(	22658	)	,
(	22669	)	,
(	22679	)	,
(	22690	)	,
(	22701	)	,
(	22712	)	,
(	22723	)	,
(	22734	)	,
(	22744	)	,
(	22755	)	,
(	22766	)	,
(	22777	)	,
(	22788	)	,
(	22799	)	,
(	22810	)	,
(	22821	)	,
(	22832	)	,
(	22843	)	,
(	22853	)	,
(	22864	)	,
(	22875	)	,
(	22886	)	,
(	22897	)	,
(	22908	)	,
(	22919	)	,
(	22930	)	,
(	22941	)	,
(	22952	)	,
(	22963	)	,
(	22974	)	,
(	22985	)	,
(	22996	)	,
(	23007	)	,
(	23018	)	,
(	23029	)	,
(	23040	)	,
(	23051	)	,
(	23062	)	,
(	23073	)	,
(	23084	)	,
(	23095	)	,
(	23106	)	,
(	23117	)	,
(	23128	)	,
(	23139	)	,
(	23150	)	,
(	23161	)	,
(	23173	)	,
(	23184	)	,
(	23195	)	,
(	23206	)	,
(	23217	)	,
(	23228	)	,
(	23239	)	,
(	23250	)	,
(	23261	)	,
(	23272	)	,
(	23284	)	,
(	23295	)	,
(	23306	)	,
(	23317	)	,
(	23328	)	,
(	23339	)	,
(	23350	)	,
(	23362	)	,
(	23373	)	,
(	23384	)	,
(	23395	)	,
(	23406	)	,
(	23417	)	,
(	23429	)	,
(	23440	)	,
(	23451	)	,
(	23462	)	,
(	23474	)	,
(	23485	)	,
(	23496	)	,
(	23507	)	,
(	23518	)	,
(	23530	)	,
(	23541	)	,
(	23552	)	,
(	23563	)	,
(	23575	)	,
(	23586	)	,
(	23597	)	,
(	23609	)	,
(	23620	)	,
(	23631	)	,
(	23642	)	,
(	23654	)	,
(	23665	)	,
(	23676	)	,
(	23688	)	,
(	23699	)	,
(	23710	)	,
(	23722	)	,
(	23733	)	,
(	23744	)	,
(	23756	)	,
(	23767	)	,
(	23778	)	,
(	23790	)	,
(	23801	)	,
(	23813	)	,
(	23824	)	,
(	23835	)	,
(	23847	)	,
(	23858	)	,
(	23870	)	,
(	23881	)	,
(	23892	)	,
(	23904	)	,
(	23915	)	,
(	23927	)	,
(	23938	)	,
(	23950	)	,
(	23961	)	,
(	23972	)	,
(	23984	)	,
(	23995	)	,
(	24007	)	,
(	24018	)	,
(	24030	)	,
(	24041	)	,
(	24053	)	,
(	24064	)	,
(	24076	)	,
(	24087	)	,
(	24099	)	,
(	24110	)	,
(	24122	)	,
(	24133	)	,
(	24145	)	,
(	24157	)	,
(	24168	)	,
(	24180	)	,
(	24191	)	,
(	24203	)	,
(	24214	)	,
(	24226	)	,
(	24238	)	,
(	24249	)	,
(	24261	)	,
(	24272	)	,
(	24284	)	,
(	24296	)	,
(	24307	)	,
(	24319	)	,
(	24330	)	,
(	24342	)	,
(	24354	)	,
(	24365	)	,
(	24377	)	,
(	24389	)	,
(	24400	)	,
(	24412	)	,
(	24424	)	,
(	24435	)	,
(	24447	)	,
(	24459	)	,
(	24470	)	,
(	24482	)	,
(	24494	)	,
(	24505	)	,
(	24517	)	,
(	24529	)	,
(	24541	)	,
(	24552	)	,
(	24564	)	,
(	24576	)	,
(	24588	)	,
(	24599	)	,
(	24611	)	,
(	24623	)	,
(	24635	)	,
(	24646	)	,
(	24658	)	,
(	24670	)	,
(	24682	)	,
(	24694	)	,
(	24705	)	,
(	24717	)	,
(	24729	)	,
(	24741	)	,
(	24753	)	,
(	24765	)	,
(	24776	)	,
(	24788	)	,
(	24800	)	,
(	24812	)	,
(	24824	)	,
(	24836	)	,
(	24848	)	,
(	24859	)	,
(	24871	)	,
(	24883	)	,
(	24895	)	,
(	24907	)	,
(	24919	)	,
(	24931	)	,
(	24943	)	,
(	24955	)	,
(	24967	)	,
(	24979	)	,
(	24990	)	,
(	25002	)	,
(	25014	)	,
(	25026	)	,
(	25038	)	,
(	25050	)	,
(	25062	)	,
(	25074	)	,
(	25086	)	,
(	25098	)	,
(	25110	)	,
(	25122	)	,
(	25134	)	,
(	25146	)	,
(	25158	)	,
(	25170	)	,
(	25182	)	,
(	25194	)	,
(	25206	)	,
(	25219	)	,
(	25231	)	,
(	25243	)	,
(	25255	)	,
(	25267	)	,
(	25279	)	,
(	25291	)	,
(	25303	)	,
(	25315	)	,
(	25327	)	,
(	25339	)	,
(	25351	)	,
(	25364	)	,
(	25376	)	,
(	25388	)	,
(	25400	)	,
(	25412	)	,
(	25424	)	,
(	25436	)	,
(	25449	)	,
(	25461	)	,
(	25473	)	,
(	25485	)	,
(	25497	)	,
(	25509	)	,
(	25522	)	,
(	25534	)	,
(	25546	)	,
(	25558	)	,
(	25571	)	,
(	25583	)	,
(	25595	)	,
(	25607	)	,
(	25619	)	,
(	25632	)	,
(	25644	)	,
(	25656	)	,
(	25669	)	,
(	25681	)	,
(	25693	)	,
(	25705	)	,
(	25718	)	,
(	25730	)	,
(	25742	)	,
(	25755	)	,
(	25767	)	,
(	25779	)	,
(	25792	)	,
(	25804	)	,
(	25816	)	,
(	25829	)	,
(	25841	)	,
(	25853	)	,
(	25866	)	,
(	25878	)	,
(	25890	)	,
(	25903	)	,
(	25915	)	,
(	25927	)	,
(	25940	)	,
(	25952	)	,
(	25965	)	,
(	25977	)	,
(	25990	)	,
(	26002	)	,
(	26014	)	,
(	26027	)	,
(	26039	)	,
(	26052	)	,
(	26064	)	,
(	26077	)	,
(	26089	)	,
(	26102	)	,
(	26114	)	,
(	26127	)	,
(	26139	)	,
(	26152	)	,
(	26164	)	,
(	26177	)	,
(	26189	)	,
(	26202	)	,
(	26214	)	,
(	26227	)	,
(	26239	)	,
(	26252	)	,
(	26264	)	,
(	26277	)	,
(	26289	)	,
(	26302	)	,
(	26315	)	,
(	26327	)	,
(	26340	)	,
(	26352	)	,
(	26365	)	,
(	26378	)	,
(	26390	)	,
(	26403	)	,
(	26415	)	,
(	26428	)	,
(	26441	)	,
(	26453	)	,
(	26466	)	,
(	26479	)	,
(	26491	)	,
(	26504	)	,
(	26517	)	,
(	26529	)	,
(	26542	)	,
(	26555	)	,
(	26567	)	,
(	26580	)	,
(	26593	)	,
(	26605	)	,
(	26618	)	,
(	26631	)	,
(	26644	)	,
(	26656	)	,
(	26669	)	,
(	26682	)	,
(	26695	)	,
(	26707	)	,
(	26720	)	,
(	26733	)	,
(	26746	)	,
(	26759	)	,
(	26771	)	,
(	26784	)	,
(	26797	)	,
(	26810	)	,
(	26823	)	,
(	26835	)	,
(	26848	)	,
(	26861	)	,
(	26874	)	,
(	26887	)	,
(	26900	)	,
(	26912	)	,
(	26925	)	,
(	26938	)	,
(	26951	)	,
(	26964	)	,
(	26977	)	,
(	26990	)	,
(	27003	)	,
(	27016	)	,
(	27029	)	,
(	27041	)	,
(	27054	)	,
(	27067	)	,
(	27080	)	,
(	27093	)	,
(	27106	)	,
(	27119	)	,
(	27132	)	,
(	27145	)	,
(	27158	)	,
(	27171	)	,
(	27184	)	,
(	27197	)	,
(	27210	)	,
(	27223	)	,
(	27236	)	,
(	27249	)	,
(	27262	)	,
(	27275	)	,
(	27288	)	,
(	27301	)	,
(	27314	)	,
(	27327	)	,
(	27340	)	,
(	27353	)	,
(	27367	)	,
(	27380	)	,
(	27393	)	,
(	27406	)	,
(	27419	)	,
(	27432	)	,
(	27445	)	,
(	27458	)	,
(	27471	)	,
(	27485	)	,
(	27498	)	,
(	27511	)	,
(	27524	)	,
(	27537	)	,
(	27550	)	,
(	27563	)	,
(	27577	)	,
(	27590	)	,
(	27603	)	,
(	27616	)	,
(	27629	)	,
(	27643	)	,
(	27656	)	,
(	27669	)	,
(	27682	)	,
(	27696	)	,
(	27709	)	,
(	27722	)	,
(	27735	)	,
(	27749	)	,
(	27762	)	,
(	27775	)	,
(	27788	)	,
(	27802	)	,
(	27815	)	,
(	27828	)	,
(	27842	)	,
(	27855	)	,
(	27868	)	,
(	27882	)	,
(	27895	)	,
(	27908	)	,
(	27922	)	,
(	27935	)	,
(	27948	)	,
(	27962	)	,
(	27975	)	,
(	27988	)	,
(	28002	)	,
(	28015	)	,
(	28029	)	,
(	28042	)	,
(	28055	)	,
(	28069	)	,
(	28082	)	,
(	28096	)	,
(	28109	)	,
(	28122	)	,
(	28136	)	,
(	28149	)	,
(	28163	)	,
(	28176	)	,
(	28190	)	,
(	28203	)	,
(	28217	)	,
(	28230	)	,
(	28244	)	,
(	28257	)	,
(	28271	)	,
(	28284	)	,
(	28298	)	,
(	28311	)	,
(	28325	)	,
(	28338	)	,
(	28352	)	,
(	28366	)	,
(	28379	)	,
(	28393	)	,
(	28406	)	,
(	28420	)	,
(	28433	)	,
(	28447	)	,
(	28461	)	,
(	28474	)	,
(	28488	)	,
(	28501	)	,
(	28515	)	,
(	28529	)	,
(	28542	)	,
(	28556	)	,
(	28570	)	,
(	28583	)	,
(	28597	)	,
(	28611	)	,
(	28624	)	,
(	28638	)	,
(	28652	)	,
(	28665	)	,
(	28679	)	,
(	28693	)	,
(	28707	)	,
(	28720	)	,
(	28734	)	,
(	28748	)	,
(	28761	)	,
(	28775	)	,
(	28789	)	,
(	28803	)	,
(	28817	)	,
(	28830	)	,
(	28844	)	,
(	28858	)	,
(	28872	)	,
(	28885	)	,
(	28899	)	,
(	28913	)	,
(	28927	)	,
(	28941	)	,
(	28955	)	,
(	28968	)	,
(	28982	)	,
(	28996	)	,
(	29010	)	,
(	29024	)	,
(	29038	)	,
(	29052	)	,
(	29066	)	,
(	29079	)	,
(	29093	)	,
(	29107	)	,
(	29121	)	,
(	29135	)	,
(	29149	)	,
(	29163	)	,
(	29177	)	,
(	29191	)	,
(	29205	)	,
(	29219	)	,
(	29233	)	,
(	29247	)	,
(	29261	)	,
(	29275	)	,
(	29289	)	,
(	29303	)	,
(	29317	)	,
(	29331	)	,
(	29345	)	,
(	29359	)	,
(	29373	)	,
(	29387	)	,
(	29401	)	,
(	29415	)	,
(	29429	)	,
(	29443	)	,
(	29457	)	,
(	29471	)	,
(	29485	)	,
(	29499	)	,
(	29514	)	,
(	29528	)	,
(	29542	)	,
(	29556	)	,
(	29570	)	,
(	29584	)	,
(	29598	)	,
(	29613	)	,
(	29627	)	,
(	29641	)	,
(	29655	)	,
(	29669	)	,
(	29683	)	,
(	29698	)	,
(	29712	)	,
(	29726	)	,
(	29740	)	,
(	29754	)	,
(	29769	)	,
(	29783	)	,
(	29797	)	,
(	29811	)	,
(	29826	)	,
(	29840	)	,
(	29854	)	,
(	29868	)	,
(	29883	)	,
(	29897	)	,
(	29911	)	,
(	29926	)	,
(	29940	)	,
(	29954	)	,
(	29969	)	,
(	29983	)	,
(	29997	)	,
(	30012	)	,
(	30026	)	,
(	30040	)	,
(	30055	)	,
(	30069	)	,
(	30083	)	,
(	30098	)	,
(	30112	)	,
(	30127	)	,
(	30141	)	,
(	30155	)	,
(	30170	)	,
(	30184	)	,
(	30199	)	,
(	30213	)	,
(	30228	)	,
(	30242	)	,
(	30256	)	,
(	30271	)	,
(	30285	)	,
(	30300	)	,
(	30314	)	,
(	30329	)	,
(	30343	)	,
(	30358	)	,
(	30372	)	,
(	30387	)	,
(	30401	)	,
(	30416	)	,
(	30430	)	,
(	30445	)	,
(	30460	)	,
(	30474	)	,
(	30489	)	,
(	30503	)	,
(	30518	)	,
(	30532	)	,
(	30547	)	,
(	30562	)	,
(	30576	)	,
(	30591	)	,
(	30606	)	,
(	30620	)	,
(	30635	)	,
(	30649	)	,
(	30664	)	,
(	30679	)	,
(	30693	)	,
(	30708	)	,
(	30723	)	,
(	30738	)	,
(	30752	)	,
(	30767	)	,
(	30782	)	,
(	30796	)	,
(	30811	)	,
(	30826	)	,
(	30841	)	,
(	30855	)	,
(	30870	)	,
(	30885	)	,
(	30900	)	,
(	30914	)	,
(	30929	)	,
(	30944	)	,
(	30959	)	,
(	30974	)	,
(	30988	)	,
(	31003	)	,
(	31018	)	,
(	31033	)	,
(	31048	)	,
(	31062	)	,
(	31077	)	,
(	31092	)	,
(	31107	)	,
(	31122	)	,
(	31137	)	,
(	31152	)	,
(	31167	)	,
(	31181	)	,
(	31196	)	,
(	31211	)	,
(	31226	)	,
(	31241	)	,
(	31256	)	,
(	31271	)	,
(	31286	)	,
(	31301	)	,
(	31316	)	,
(	31331	)	,
(	31346	)	,
(	31361	)	,
(	31376	)	,
(	31391	)	,
(	31406	)	,
(	31421	)	,
(	31436	)	,
(	31451	)	,
(	31466	)	,
(	31481	)	,
(	31496	)	,
(	31511	)	,
(	31526	)	,
(	31541	)	,
(	31556	)	,
(	31571	)	,
(	31587	)	,
(	31602	)	,
(	31617	)	,
(	31632	)	,
(	31647	)	,
(	31662	)	,
(	31677	)	,
(	31692	)	,
(	31708	)	,
(	31723	)	,
(	31738	)	,
(	31753	)	,
(	31768	)	,
(	31783	)	,
(	31799	)	,
(	31814	)	,
(	31829	)	,
(	31844	)	,
(	31860	)	,
(	31875	)	,
(	31890	)	,
(	31905	)	,
(	31920	)	,
(	31936	)	,
(	31951	)	,
(	31966	)	,
(	31982	)	,
(	31997	)	,
(	32012	)	,
(	32027	)	,
(	32043	)	,
(	32058	)	,
(	32073	)	,
(	32089	)	,
(	32104	)	,
(	32119	)	,
(	32135	)	,
(	32150	)	,
(	32166	)	,
(	32181	)	,
(	32196	)	,
(	32212	)	,
(	32227	)	,
(	32243	)	,
(	32258	)	,
(	32273	)	,
(	32289	)	,
(	32304	)	,
(	32320	)	,
(	32335	)	,
(	32351	)	,
(	32366	)	,
(	32382	)	,
(	32397	)	,
(	32413	)	,
(	32428	)	,
(	32444	)	,
(	32459	)	,
(	32475	)	,
(	32490	)	,
(	32506	)	,
(	32521	)	,
(	32537	)	,
(	32552	)	,
(	32568	)	,
(	32583	)	,
(	32599	)	,
(	32615	)	,
(	32630	)	,
(	32646	)	,
(	32661	)	,
(	32677	)	,
(	32693	)	,
(	32708	)	,
(	32724	)	,
(	32740	)	,
(	32755	)	,
(	32771	)	,
(	32787	)	,
(	32802	)	,
(	32818	)	,
(	32834	)	,
(	32849	)	,
(	32865	)	,
(	32881	)	,
(	32896	)	,
(	32912	)	,
(	32928	)	,
(	32944	)	,
(	32959	)	,
(	32975	)	,
(	32991	)	,
(	33007	)	,
(	33022	)	,
(	33038	)	,
(	33054	)	,
(	33070	)	,
(	33086	)	,
(	33101	)	,
(	33117	)	,
(	33133	)	,
(	33149	)	,
(	33165	)	,
(	33181	)	,
(	33197	)	,
(	33212	)	,
(	33228	)	,
(	33244	)	,
(	33260	)	,
(	33276	)	,
(	33292	)	,
(	33308	)	,
(	33324	)	,
(	33340	)	,
(	33356	)	,
(	33372	)	,
(	33388	)	,
(	33404	)	,
(	33419	)	,
(	33435	)	,
(	33451	)	,
(	33467	)	,
(	33483	)	,
(	33499	)	,
(	33515	)	,
(	33532	)	,
(	33548	)	,
(	33564	)	,
(	33580	)	,
(	33596	)	,
(	33612	)	,
(	33628	)	,
(	33644	)	,
(	33660	)	,
(	33676	)	,
(	33692	)	,
(	33708	)	,
(	33724	)	,
(	33741	)	,
(	33757	)	,
(	33773	)	,
(	33789	)	,
(	33805	)	,
(	33821	)	,
(	33837	)	,
(	33854	)	,
(	33870	)	,
(	33886	)	,
(	33902	)	,
(	33918	)	,
(	33935	)	,
(	33951	)	,
(	33967	)	,
(	33983	)	,
(	34000	)	,
(	34016	)	,
(	34032	)	,
(	34048	)	,
(	34065	)	,
(	34081	)	,
(	34097	)	,
(	34114	)	,
(	34130	)	,
(	34146	)	,
(	34163	)	,
(	34179	)	,
(	34195	)	,
(	34212	)	,
(	34228	)	,
(	34244	)	,
(	34261	)	,
(	34277	)	,
(	34293	)	,
(	34310	)	,
(	34326	)	,
(	34343	)	,
(	34359	)	,
(	34375	)	,
(	34392	)	,
(	34408	)	,
(	34425	)	,
(	34441	)	,
(	34458	)	,
(	34474	)	,
(	34491	)	,
(	34507	)	,
(	34524	)	,
(	34540	)	,
(	34557	)	,
(	34573	)	,
(	34590	)	,
(	34606	)	,
(	34623	)	,
(	34639	)	,
(	34656	)	,
(	34673	)	,
(	34689	)	,
(	34706	)	,
(	34722	)	,
(	34739	)	,
(	34756	)	,
(	34772	)	,
(	34789	)	,
(	34805	)	,
(	34822	)	,
(	34839	)	,
(	34855	)	,
(	34872	)	,
(	34889	)	,
(	34905	)	,
(	34922	)	,
(	34939	)	,
(	34955	)	,
(	34972	)	,
(	34989	)	,
(	35006	)	,
(	35022	)	,
(	35039	)	,
(	35056	)	,
(	35073	)	,
(	35089	)	,
(	35106	)	,
(	35123	)	,
(	35140	)	,
(	35157	)	,
(	35173	)	,
(	35190	)	,
(	35207	)	,
(	35224	)	,
(	35241	)	,
(	35258	)	,
(	35274	)	,
(	35291	)	,
(	35308	)	,
(	35325	)	,
(	35342	)	,
(	35359	)	,
(	35376	)	,
(	35393	)	,
(	35410	)	,
(	35426	)	,
(	35443	)	,
(	35460	)	,
(	35477	)	,
(	35494	)	,
(	35511	)	,
(	35528	)	,
(	35545	)	,
(	35562	)	,
(	35579	)	,
(	35596	)	,
(	35613	)	,
(	35630	)	,
(	35647	)	,
(	35664	)	,
(	35681	)	,
(	35698	)	,
(	35716	)	,
(	35733	)	,
(	35750	)	,
(	35767	)	,
(	35784	)	,
(	35801	)	,
(	35818	)	,
(	35835	)	,
(	35852	)	,
(	35870	)	,
(	35887	)	,
(	35904	)	,
(	35921	)	,
(	35938	)	,
(	35955	)	,
(	35973	)	,
(	35990	)	,
(	36007	)	,
(	36024	)	,
(	36041	)	,
(	36059	)	,
(	36076	)	,
(	36093	)	,
(	36110	)	,
(	36128	)	,
(	36145	)	,
(	36162	)	,
(	36179	)	,
(	36197	)	,
(	36214	)	,
(	36231	)	,
(	36249	)	,
(	36266	)	,
(	36283	)	,
(	36301	)	,
(	36318	)	,
(	36335	)	,
(	36353	)	,
(	36370	)	,
(	36388	)	,
(	36405	)	,
(	36422	)	,
(	36440	)	,
(	36457	)	,
(	36475	)	,
(	36492	)	,
(	36510	)	,
(	36527	)	,
(	36545	)	,
(	36562	)	,
(	36579	)	,
(	36597	)	,
(	36614	)	,
(	36632	)	,
(	36649	)	,
(	36667	)	,
(	36685	)	,
(	36702	)	,
(	36720	)	,
(	36737	)	,
(	36755	)	,
(	36772	)	,
(	36790	)	,
(	36808	)	,
(	36825	)	,
(	36843	)	,
(	36860	)	,
(	36878	)	,
(	36896	)	,
(	36913	)	,
(	36931	)	,
(	36949	)	,
(	36966	)	,
(	36984	)	,
(	37002	)	,
(	37019	)	,
(	37037	)	,
(	37055	)	,
(	37072	)	,
(	37090	)	,
(	37108	)	,
(	37126	)	,
(	37143	)	,
(	37161	)	,
(	37179	)	,
(	37197	)	,
(	37214	)	,
(	37232	)	,
(	37250	)	,
(	37268	)	,
(	37286	)	,
(	37303	)	,
(	37321	)	,
(	37339	)	,
(	37357	)	,
(	37375	)	,
(	37393	)	,
(	37411	)	,
(	37429	)	,
(	37446	)	,
(	37464	)	,
(	37482	)	,
(	37500	)	,
(	37518	)	,
(	37536	)	,
(	37554	)	,
(	37572	)	,
(	37590	)	,
(	37608	)	,
(	37626	)	,
(	37644	)	,
(	37662	)	,
(	37680	)	,
(	37698	)	,
(	37716	)	,
(	37734	)	,
(	37752	)	,
(	37770	)	,
(	37788	)	,
(	37806	)	,
(	37824	)	,
(	37842	)	,
(	37860	)	,
(	37879	)	,
(	37897	)	,
(	37915	)	,
(	37933	)	,
(	37951	)	,
(	37969	)	,
(	37987	)	,
(	38005	)	,
(	38024	)	,
(	38042	)	,
(	38060	)	,
(	38078	)	,
(	38096	)	,
(	38115	)	,
(	38133	)	,
(	38151	)	,
(	38169	)	,
(	38188	)	,
(	38206	)	,
(	38224	)	,
(	38242	)	,
(	38261	)	,
(	38279	)	,
(	38297	)	,
(	38316	)	,
(	38334	)	,
(	38352	)	,
(	38371	)	,
(	38389	)	,
(	38407	)	,
(	38426	)	,
(	38444	)	,
(	38462	)	,
(	38481	)	,
(	38499	)	,
(	38518	)	,
(	38536	)	,
(	38554	)	,
(	38573	)	,
(	38591	)	,
(	38610	)	,
(	38628	)	,
(	38647	)	,
(	38665	)	,
(	38684	)	,
(	38702	)	,
(	38721	)	,
(	38739	)	,
(	38758	)	,
(	38776	)	,
(	38795	)	,
(	38813	)	,
(	38832	)	,
(	38850	)	,
(	38869	)	,
(	38888	)	,
(	38906	)	,
(	38925	)	,
(	38943	)	,
(	38962	)	,
(	38981	)	,
(	38999	)	,
(	39018	)	,
(	39037	)	,
(	39055	)	,
(	39074	)	,
(	39093	)	,
(	39111	)	,
(	39130	)	,
(	39149	)	,
(	39167	)	,
(	39186	)	,
(	39205	)	,
(	39224	)	,
(	39242	)	,
(	39261	)	,
(	39280	)	,
(	39299	)	,
(	39318	)	,
(	39336	)	,
(	39355	)	,
(	39374	)	,
(	39393	)	,
(	39412	)	,
(	39430	)	,
(	39449	)	,
(	39468	)	,
(	39487	)	,
(	39506	)	,
(	39525	)	,
(	39544	)	,
(	39563	)	,
(	39582	)	,
(	39600	)	,
(	39619	)	,
(	39638	)	,
(	39657	)	,
(	39676	)	,
(	39695	)	,
(	39714	)	,
(	39733	)	,
(	39752	)	,
(	39771	)	,
(	39790	)	,
(	39809	)	,
(	39828	)	,
(	39847	)	,
(	39866	)	,
(	39885	)	,
(	39905	)	,
(	39924	)	,
(	39943	)	,
(	39962	)	,
(	39981	)	,
(	40000	)	,
(	40019	)	,
(	40038	)	,
(	40057	)	,
(	40077	)	,
(	40096	)	,
(	40115	)	,
(	40134	)	,
(	40153	)	,
(	40172	)	,
(	40192	)	,
(	40211	)	,
(	40230	)	,
(	40249	)	,
(	40269	)	,
(	40288	)	,
(	40307	)	,
(	40326	)	,
(	40346	)	,
(	40365	)	,
(	40384	)	,
(	40404	)	,
(	40423	)	,
(	40442	)	,
(	40462	)	,
(	40481	)	,
(	40500	)	,
(	40520	)	,
(	40539	)	,
(	40558	)	,
(	40578	)	,
(	40597	)	,
(	40617	)	,
(	40636	)	,
(	40655	)	,
(	40675	)	,
(	40694	)	,
(	40714	)	,
(	40733	)	,
(	40753	)	,
(	40772	)	,
(	40792	)	,
(	40811	)	,
(	40831	)	,
(	40850	)	,
(	40870	)	,
(	40889	)	,
(	40909	)	,
(	40928	)	,
(	40948	)	,
(	40968	)	,
(	40987	)	,
(	41007	)	,
(	41026	)	,
(	41046	)	,
(	41066	)	,
(	41085	)	,
(	41105	)	,
(	41125	)	,
(	41144	)	,
(	41164	)	,
(	41184	)	,
(	41203	)	,
(	41223	)	,
(	41243	)	,
(	41262	)	,
(	41282	)	,
(	41302	)	,
(	41322	)	,
(	41341	)	,
(	41361	)	,
(	41381	)	,
(	41401	)	,
(	41420	)	,
(	41440	)	,
(	41460	)	,
(	41480	)	,
(	41500	)	,
(	41520	)	,
(	41539	)	,
(	41559	)	,
(	41579	)	,
(	41599	)	,
(	41619	)	,
(	41639	)	,
(	41659	)	,
(	41679	)	,
(	41699	)	,
(	41719	)	,
(	41739	)	,
(	41758	)	,
(	41778	)	,
(	41798	)	,
(	41818	)	,
(	41838	)	,
(	41858	)	,
(	41878	)	,
(	41898	)	,
(	41918	)	,
(	41939	)	,
(	41959	)	,
(	41979	)	,
(	41999	)	,
(	42019	)	,
(	42039	)	,
(	42059	)	,
(	42079	)	,
(	42099	)	,
(	42119	)	,
(	42139	)	,
(	42160	)	,
(	42180	)	,
(	42200	)	,
(	42220	)	,
(	42240	)	,
(	42261	)	,
(	42281	)	,
(	42301	)	,
(	42321	)	,
(	42341	)	,
(	42362	)	,
(	42382	)	,
(	42402	)	,
(	42422	)	,
(	42443	)	,
(	42463	)	,
(	42483	)	,
(	42504	)	,
(	42524	)	,
(	42544	)	,
(	42565	)	,
(	42585	)	,
(	42605	)	,
(	42626	)	,
(	42646	)	,
(	42666	)	,
(	42687	)	,
(	42707	)	,
(	42728	)	,
(	42748	)	,
(	42769	)	,
(	42789	)	,
(	42810	)	,
(	42830	)	,
(	42850	)	,
(	42871	)	,
(	42891	)	,
(	42912	)	,
(	42932	)	,
(	42953	)	,
(	42974	)	,
(	42994	)	,
(	43015	)	,
(	43035	)	,
(	43056	)	,
(	43076	)	,
(	43097	)	,
(	43118	)	,
(	43138	)	,
(	43159	)	,
(	43179	)	,
(	43200	)	,
(	43221	)	,
(	43241	)	,
(	43262	)	,
(	43283	)	,
(	43303	)	,
(	43324	)	,
(	43345	)	,
(	43366	)	,
(	43386	)	,
(	43407	)	,
(	43428	)	,
(	43449	)	,
(	43469	)	,
(	43490	)	,
(	43511	)	,
(	43532	)	,
(	43553	)	,
(	43573	)	,
(	43594	)	,
(	43615	)	,
(	43636	)	,
(	43657	)	,
(	43678	)	,
(	43699	)	,
(	43719	)	,
(	43740	)	,
(	43761	)	,
(	43782	)	,
(	43803	)	,
(	43824	)	,
(	43845	)	,
(	43866	)	,
(	43887	)	,
(	43908	)	,
(	43929	)	,
(	43950	)	,
(	43971	)	,
(	43992	)	,
(	44013	)	,
(	44034	)	,
(	44055	)	,
(	44076	)	,
(	44097	)	,
(	44118	)	,
(	44139	)	,
(	44161	)	,
(	44182	)	,
(	44203	)	,
(	44224	)	,
(	44245	)	,
(	44266	)	,
(	44287	)	,
(	44309	)	,
(	44330	)	,
(	44351	)	,
(	44372	)	,
(	44393	)	,
(	44415	)	,
(	44436	)	,
(	44457	)	,
(	44478	)	,
(	44500	)	,
(	44521	)	,
(	44542	)	,
(	44563	)	,
(	44585	)	,
(	44606	)	,
(	44627	)	,
(	44649	)	,
(	44670	)	,
(	44691	)	,
(	44713	)	,
(	44734	)	,
(	44756	)	,
(	44777	)	,
(	44798	)	,
(	44820	)	,
(	44841	)	,
(	44863	)	,
(	44884	)	,
(	44906	)	,
(	44927	)	,
(	44949	)	,
(	44970	)	,
(	44992	)	,
(	45013	)	,
(	45035	)	,
(	45056	)	,
(	45078	)	,
(	45099	)	,
(	45121	)	,
(	45142	)	,
(	45164	)	,
(	45186	)	,
(	45207	)	,
(	45229	)	,
(	45250	)	,
(	45272	)	,
(	45294	)	,
(	45315	)	,
(	45337	)	,
(	45359	)	,
(	45380	)	,
(	45402	)	,
(	45424	)	,
(	45446	)	,
(	45467	)	,
(	45489	)	,
(	45511	)	,
(	45532	)	,
(	45554	)	,
(	45576	)	,
(	45598	)	,
(	45620	)	,
(	45641	)	,
(	45663	)	,
(	45685	)	,
(	45707	)	,
(	45729	)	,
(	45751	)	,
(	45773	)	,
(	45794	)	,
(	45816	)	,
(	45838	)	,
(	45860	)	,
(	45882	)	,
(	45904	)	,
(	45926	)	,
(	45948	)	,
(	45970	)	,
(	45992	)	,
(	46014	)	,
(	46036	)	,
(	46058	)	,
(	46080	)	,
(	46102	)	,
(	46124	)	,
(	46146	)	,
(	46168	)	,
(	46190	)	,
(	46212	)	,
(	46234	)	,
(	46256	)	,
(	46279	)	,
(	46301	)	,
(	46323	)	,
(	46345	)	,
(	46367	)	,
(	46389	)	,
(	46412	)	,
(	46434	)	,
(	46456	)	,
(	46478	)	,
(	46500	)	,
(	46523	)	,
(	46545	)	,
(	46567	)	,
(	46589	)	,
(	46612	)	,
(	46634	)	,
(	46656	)	,
(	46679	)	,
(	46701	)	,
(	46723	)	,
(	46746	)	,
(	46768	)	,
(	46790	)	,
(	46813	)	,
(	46835	)	,
(	46857	)	,
(	46880	)	,
(	46902	)	,
(	46925	)	,
(	46947	)	,
(	46969	)	,
(	46992	)	,
(	47014	)	,
(	47037	)	,
(	47059	)	,
(	47082	)	,
(	47104	)	,
(	47127	)	,
(	47149	)	,
(	47172	)	,
(	47195	)	,
(	47217	)	,
(	47240	)	,
(	47262	)	,
(	47285	)	,
(	47308	)	,
(	47330	)	,
(	47353	)	,
(	47375	)	,
(	47398	)	,
(	47421	)	,
(	47443	)	,
(	47466	)	,
(	47489	)	,
(	47511	)	,
(	47534	)	,
(	47557	)	,
(	47580	)	,
(	47602	)	,
(	47625	)	,
(	47648	)	,
(	47671	)	,
(	47694	)	,
(	47716	)	,
(	47739	)	,
(	47762	)	,
(	47785	)	,
(	47808	)	,
(	47831	)	,
(	47853	)	,
(	47876	)	,
(	47899	)	,
(	47922	)	,
(	47945	)	,
(	47968	)	,
(	47991	)	,
(	48014	)	,
(	48037	)	,
(	48060	)	,
(	48083	)	,
(	48106	)	,
(	48129	)	,
(	48152	)	,
(	48175	)	,
(	48198	)	,
(	48221	)	,
(	48244	)	,
(	48267	)	,
(	48290	)	,
(	48313	)	,
(	48336	)	,
(	48359	)	,
(	48382	)	,
(	48406	)	,
(	48429	)	,
(	48452	)	,
(	48475	)	,
(	48498	)	,
(	48521	)	,
(	48545	)	,
(	48568	)	,
(	48591	)	,
(	48614	)	,
(	48637	)	,
(	48661	)	,
(	48684	)	,
(	48707	)	,
(	48731	)	,
(	48754	)	,
(	48777	)	,
(	48801	)	,
(	48824	)	,
(	48847	)	,
(	48871	)	,
(	48894	)	,
(	48917	)	,
(	48941	)	,
(	48964	)	,
(	48988	)	,
(	49011	)	,
(	49034	)	,
(	49058	)	,
(	49081	)	,
(	49105	)	,
(	49128	)	,
(	49152	)	,
(	49175	)	,
(	49199	)	,
(	49222	)	,
(	49246	)	,
(	49269	)	,
(	49293	)	,
(	49316	)	,
(	49340	)	,
(	49364	)	,
(	49387	)	,
(	49411	)	,
(	49434	)	,
(	49458	)	,
(	49482	)	,
(	49505	)	,
(	49529	)	,
(	49553	)	,
(	49576	)	,
(	49600	)	,
(	49624	)	,
(	49648	)	,
(	49671	)	,
(	49695	)	,
(	49719	)	,
(	49743	)	,
(	49766	)	,
(	49790	)	,
(	49814	)	,
(	49838	)	,
(	49862	)	,
(	49886	)	,
(	49909	)	,
(	49933	)	,
(	49957	)	,
(	49981	)	,
(	50005	)	,
(	50029	)	,
(	50053	)	,
(	50077	)	,
(	50101	)	,
(	50125	)	,
(	50149	)	,
(	50172	)	,
(	50196	)	,
(	50220	)	,
(	50244	)	,
(	50269	)	,
(	50293	)	,
(	50317	)	,
(	50341	)	,
(	50365	)	,
(	50389	)	,
(	50413	)	,
(	50437	)	,
(	50461	)	,
(	50485	)	,
(	50509	)	,
(	50534	)	,
(	50558	)	,
(	50582	)	,
(	50606	)	,
(	50630	)	,
(	50654	)	,
(	50679	)	,
(	50703	)	,
(	50727	)	,
(	50751	)	,
(	50776	)	,
(	50800	)	,
(	50824	)	,
(	50849	)	,
(	50873	)	,
(	50897	)	,
(	50922	)	,
(	50946	)	,
(	50970	)	,
(	50995	)	,
(	51019	)	,
(	51043	)	,
(	51068	)	,
(	51092	)	,
(	51117	)	,
(	51141	)	,
(	51166	)	,
(	51190	)	,
(	51214	)	,
(	51239	)	,
(	51263	)	,
(	51288	)	,
(	51313	)	,
(	51337	)	,
(	51362	)	,
(	51386	)	,
(	51411	)	,
(	51435	)	,
(	51460	)	,
(	51484	)	,
(	51509	)	,
(	51534	)	,
(	51558	)	,
(	51583	)	,
(	51608	)	,
(	51632	)	,
(	51657	)	,
(	51682	)	,
(	51706	)	,
(	51731	)	,
(	51756	)	,
(	51781	)	,
(	51805	)	,
(	51830	)	,
(	51855	)	,
(	51880	)	,
(	51905	)	,
(	51929	)	,
(	51954	)	,
(	51979	)	,
(	52004	)	,
(	52029	)	,
(	52054	)	,
(	52079	)	,
(	52103	)	,
(	52128	)	,
(	52153	)	,
(	52178	)	,
(	52203	)	,
(	52228	)	,
(	52253	)	,
(	52278	)	,
(	52303	)	,
(	52328	)	,
(	52353	)	,
(	52378	)	,
(	52403	)	,
(	52428	)	,
(	52453	)	,
(	52478	)	,
(	52504	)	,
(	52529	)	,
(	52554	)	,
(	52579	)	,
(	52604	)	,
(	52629	)	,
(	52654	)	,
(	52679	)	,
(	52705	)	,
(	52730	)	,
(	52755	)	,
(	52780	)	,
(	52806	)	,
(	52831	)	,
(	52856	)	,
(	52881	)	,
(	52907	)	,
(	52932	)	,
(	52957	)	,
(	52983	)	,
(	53008	)	,
(	53033	)	,
(	53059	)	,
(	53084	)	,
(	53109	)	,
(	53135	)	,
(	53160	)	,
(	53186	)	,
(	53211	)	,
(	53236	)	,
(	53262	)	,
(	53287	)	,
(	53313	)	,
(	53338	)	,
(	53364	)	,
(	53389	)	,
(	53415	)	,
(	53440	)	,
(	53466	)	,
(	53492	)	,
(	53517	)	,
(	53543	)	,
(	53568	)	,
(	53594	)	,
(	53620	)	,
(	53645	)	,
(	53671	)	,
(	53696	)	,
(	53722	)	,
(	53748	)	,
(	53774	)	,
(	53799	)	,
(	53825	)	,
(	53851	)	,
(	53876	)	,
(	53902	)	,
(	53928	)	,
(	53954	)	,
(	53980	)	,
(	54005	)	,
(	54031	)	,
(	54057	)	,
(	54083	)	,
(	54109	)	,
(	54135	)	,
(	54161	)	,
(	54186	)	,
(	54212	)	,
(	54238	)	,
(	54264	)	,
(	54290	)	,
(	54316	)	,
(	54342	)	,
(	54368	)	,
(	54394	)	,
(	54420	)	,
(	54446	)	,
(	54472	)	,
(	54498	)	,
(	54524	)	,
(	54550	)	,
(	54576	)	,
(	54602	)	,
(	54629	)	,
(	54655	)	,
(	54681	)	,
(	54707	)	,
(	54733	)	,
(	54759	)	,
(	54785	)	,
(	54812	)	,
(	54838	)	,
(	54864	)	,
(	54890	)	,
(	54917	)	,
(	54943	)	,
(	54969	)	,
(	54995	)	,
(	55022	)	,
(	55048	)	,
(	55074	)	,
(	55101	)	,
(	55127	)	,
(	55153	)	,
(	55180	)	,
(	55206	)	,
(	55232	)	,
(	55259	)	,
(	55285	)	,
(	55312	)	,
(	55338	)	,
(	55365	)	,
(	55391	)	,
(	55418	)	,
(	55444	)	,
(	55471	)	,
(	55497	)	,
(	55524	)	,
(	55550	)	,
(	55577	)	,
(	55603	)	,
(	55630	)	,
(	55657	)	,
(	55683	)	,
(	55710	)	,
(	55736	)	,
(	55763	)	,
(	55790	)	,
(	55816	)	,
(	55843	)	,
(	55870	)	,
(	55897	)	,
(	55923	)	,
(	55950	)	,
(	55977	)	,
(	56004	)	,
(	56030	)	,
(	56057	)	,
(	56084	)	,
(	56111	)	,
(	56138	)	,
(	56164	)	,
(	56191	)	,
(	56218	)	,
(	56245	)	,
(	56272	)	,
(	56299	)	,
(	56326	)	,
(	56353	)	,
(	56380	)	,
(	56407	)	,
(	56433	)	,
(	56460	)	,
(	56487	)	,
(	56514	)	,
(	56542	)	,
(	56569	)	,
(	56596	)	,
(	56623	)	,
(	56650	)	,
(	56677	)	,
(	56704	)	,
(	56731	)	,
(	56758	)	,
(	56785	)	,
(	56812	)	,
(	56840	)	,
(	56867	)	,
(	56894	)	,
(	56921	)	,
(	56948	)	,
(	56976	)	,
(	57003	)	,
(	57030	)	,
(	57057	)	,
(	57085	)	,
(	57112	)	,
(	57139	)	,
(	57167	)	,
(	57194	)	,
(	57221	)	,
(	57249	)	,
(	57276	)	,
(	57303	)	,
(	57331	)	,
(	57358	)	,
(	57386	)	,
(	57413	)	,
(	57441	)	,
(	57468	)	,
(	57495	)	,
(	57523	)	,
(	57550	)	,
(	57578	)	,
(	57606	)	,
(	57633	)	,
(	57661	)	,
(	57688	)	,
(	57716	)	,
(	57743	)	,
(	57771	)	,
(	57799	)	,
(	57826	)	,
(	57854	)	,
(	57882	)	,
(	57909	)	,
(	57937	)	,
(	57965	)	,
(	57992	)	,
(	58020	)	,
(	58048	)	,
(	58076	)	,
(	58103	)	,
(	58131	)	,
(	58159	)	,
(	58187	)	,
(	58215	)	,
(	58242	)	,
(	58270	)	,
(	58298	)	,
(	58326	)	,
(	58354	)	,
(	58382	)	,
(	58410	)	,
(	58438	)	,
(	58466	)	,
(	58493	)	,
(	58521	)	,
(	58549	)	,
(	58577	)	,
(	58605	)	,
(	58633	)	,
(	58661	)	,
(	58690	)	,
(	58718	)	,
(	58746	)	,
(	58774	)	,
(	58802	)	,
(	58830	)	,
(	58858	)	,
(	58886	)	,
(	58914	)	,
(	58943	)	,
(	58971	)	,
(	58999	)	,
(	59027	)	,
(	59055	)	,
(	59084	)	,
(	59112	)	,
(	59140	)	,
(	59168	)	,
(	59197	)	,
(	59225	)	,
(	59253	)	,
(	59282	)	,
(	59310	)	,
(	59338	)	,
(	59367	)	,
(	59395	)	,
(	59424	)	,
(	59452	)	,
(	59480	)	,
(	59509	)	,
(	59537	)	,
(	59566	)	,
(	59594	)	,
(	59623	)	,
(	59651	)	,
(	59680	)	,
(	59708	)	,
(	59737	)	,
(	59765	)	,
(	59794	)	,
(	59823	)	,
(	59851	)	,
(	59880	)	,
(	59908	)	,
(	59937	)	,
(	59966	)	,
(	59994	)	,
(	60023	)	,
(	60052	)	,
(	60080	)	,
(	60109	)	,
(	60138	)	,
(	60167	)	,
(	60195	)	,
(	60224	)	,
(	60253	)	,
(	60282	)	,
(	60311	)	,
(	60340	)	,
(	60368	)	,
(	60397	)	,
(	60426	)	,
(	60455	)	,
(	60484	)	,
(	60513	)	,
(	60542	)	,
(	60571	)	,
(	60600	)	,
(	60629	)	,
(	60658	)	,
(	60687	)	,
(	60716	)	,
(	60745	)	,
(	60774	)	,
(	60803	)	,
(	60832	)	,
(	60861	)	,
(	60890	)	,
(	60919	)	,
(	60948	)	,
(	60977	)	,
(	61007	)	,
(	61036	)	,
(	61065	)	,
(	61094	)	,
(	61123	)	,
(	61153	)	,
(	61182	)	,
(	61211	)	,
(	61240	)	,
(	61270	)	,
(	61299	)	,
(	61328	)	,
(	61358	)	,
(	61387	)	,
(	61416	)	,
(	61446	)	,
(	61475	)	,
(	61504	)	,
(	61534	)	,
(	61563	)	,
(	61593	)	,
(	61622	)	,
(	61652	)	,
(	61681	)	,
(	61711	)	,
(	61740	)	,
(	61770	)	,
(	61799	)	,
(	61829	)	,
(	61858	)	,
(	61888	)	,
(	61917	)	,
(	61947	)	,
(	61977	)	,
(	62006	)	,
(	62036	)	,
(	62066	)	,
(	62095	)	,
(	62125	)	,
(	62155	)	,
(	62184	)	,
(	62214	)	,
(	62244	)	,
(	62274	)	,
(	62303	)	,
(	62333	)	,
(	62363	)	,
(	62393	)	,
(	62423	)	,
(	62452	)	,
(	62482	)	,
(	62512	)	,
(	62542	)	,
(	62572	)	,
(	62602	)	,
(	62632	)	,
(	62662	)	,
(	62692	)	,
(	62722	)	,
(	62752	)	,
(	62782	)	,
(	62812	)	,
(	62842	)	,
(	62872	)	,
(	62902	)	,
(	62932	)	,
(	62962	)	,
(	62992	)	,
(	63022	)	,
(	63052	)	,
(	63083	)	,
(	63113	)	,
(	63143	)	,
(	63173	)	,
(	63203	)	,
(	63234	)	,
(	63264	)	,
(	63294	)	,
(	63324	)	,
(	63355	)	,
(	63385	)	,
(	63415	)	,
(	63445	)	,
(	63476	)	,
(	63506	)	,
(	63537	)	,
(	63567	)	,
(	63597	)	,
(	63628	)	,
(	63658	)	,
(	63689	)	,
(	63719	)	,
(	63749	)	,
(	63780	)	,
(	63810	)	,
(	63841	)	,
(	63872	)	,
(	63902	)	,
(	63933	)	,
(	63963	)	,
(	63994	)	,
(	64024	)	,
(	64055	)	,
(	64086	)	,
(	64116	)	,
(	64147	)	,
(	64178	)	,
(	64208	)	,
(	64239	)	,
(	64270	)	,
(	64300	)	,
(	64331	)	,
(	64362	)	,
(	64393	)	,
(	64423	)	,
(	64454	)	,
(	64485	)	,
(	64516	)	,
(	64547	)	,
(	64578	)	,
(	64609	)	,
(	64639	)	,
(	64670	)	,
(	64701	)	,
(	64732	)	,
(	64763	)	,
(	64794	)	,
(	64825	)	,
(	64856	)	,
(	64887	)	,
(	64918	)	,
(	64949	)	,
(	64980	)	,
(	65011	)	,
(	65042	)	,
(	65073	)	,
(	65105	)	,
(	65136	)	,
(	65167	)	,
(	65198	)	,
(	65229	)	,
(	65260	)	,
(	65292	)	,
(	65323	)	,
(	65354	)	,
(	65385	)	,
(	65417	)	,
(	65448	)	,
(	65479	)	,
(	65510	)	,
(	65542	)	,
(	65573	)	,
(	65604	)	,
(	65636	)	,
(	65667	)	,
(	65699	)	,
(	65730	)	,
(	65761	)	,
(	65793	)	,
(	65824	)	,
(	65856	)	,
(	65887	)	,
(	65919	)	,
(	65950	)	,
(	65982	)	,
(	66013	)	,
(	66045	)	,
(	66077	)	,
(	66108	)	,
(	66140	)	,
(	66171	)	,
(	66203	)	,
(	66235	)	,
(	66266	)	,
(	66298	)	,
(	66330	)	,
(	66361	)	,
(	66393	)	,
(	66425	)	,
(	66457	)	,
(	66488	)	,
(	66520	)	,
(	66552	)	,
(	66584	)	,
(	66616	)	,
(	66648	)	,
(	66679	)	,
(	66711	)	,
(	66743	)	,
(	66775	)	,
(	66807	)	,
(	66839	)	,
(	66871	)	,
(	66903	)	,
(	66935	)	,
(	66967	)	,
(	66999	)	,
(	67031	)	,
(	67063	)	,
(	67095	)	,
(	67127	)	,
(	67159	)	,
(	67191	)	,
(	67223	)	,
(	67256	)	,
(	67288	)	,
(	67320	)	,
(	67352	)	,
(	67384	)	,
(	67417	)	,
(	67449	)	,
(	67481	)	,
(	67513	)	,
(	67546	)	,
(	67578	)	,
(	67610	)	,
(	67643	)	,
(	67675	)	,
(	67707	)	,
(	67740	)	,
(	67772	)	,
(	67804	)	,
(	67837	)	,
(	67869	)	,
(	67902	)	,
(	67934	)	,
(	67967	)	,
(	67999	)	,
(	68032	)	,
(	68064	)	,
(	68097	)	,
(	68129	)	,
(	68162	)	,
(	68194	)	,
(	68227	)	,
(	68260	)	,
(	68292	)	,
(	68325	)	,
(	68358	)	,
(	68390	)	,
(	68423	)	,
(	68456	)	,
(	68489	)	,
(	68521	)	,
(	68554	)	,
(	68587	)	,
(	68620	)	,
(	68652	)	,
(	68685	)	,
(	68718	)	,
(	68751	)	,
(	68784	)	,
(	68817	)	,
(	68850	)	,
(	68883	)	,
(	68915	)	,
(	68948	)	,
(	68981	)	,
(	69014	)	,
(	69047	)	,
(	69080	)	,
(	69113	)	,
(	69146	)	,
(	69180	)	,
(	69213	)	,
(	69246	)	,
(	69279	)	,
(	69312	)	,
(	69345	)	,
(	69378	)	,
(	69411	)	,
(	69445	)	,
(	69478	)	,
(	69511	)	,
(	69544	)	,
(	69577	)	,
(	69611	)	,
(	69644	)	,
(	69677	)	,
(	69711	)	,
(	69744	)	,
(	69777	)	,
(	69811	)	,
(	69844	)	,
(	69877	)	,
(	69911	)	,
(	69944	)	,
(	69978	)	,
(	70011	)	,
(	70045	)	,
(	70078	)	,
(	70112	)	,
(	70145	)	,
(	70179	)	,
(	70212	)	,
(	70246	)	,
(	70279	)	,
(	70313	)	,
(	70347	)	,
(	70380	)	,
(	70414	)	,
(	70448	)	,
(	70481	)	,
(	70515	)	,
(	70549	)	,
(	70582	)	,
(	70616	)	,
(	70650	)	,
(	70684	)	,
(	70718	)	,
(	70751	)	,
(	70785	)	,
(	70819	)	,
(	70853	)	,
(	70887	)	,
(	70921	)	,
(	70955	)	,
(	70989	)	,
(	71022	)	,
(	71056	)	,
(	71090	)	,
(	71124	)	,
(	71158	)	,
(	71192	)	,
(	71226	)	,
(	71261	)	,
(	71295	)	,
(	71329	)	,
(	71363	)	,
(	71397	)	,
(	71431	)	,
(	71465	)	,
(	71499	)	,
(	71534	)	,
(	71568	)	,
(	71602	)	,
(	71636	)	,
(	71670	)	,
(	71705	)	,
(	71739	)	,
(	71773	)	,
(	71808	)	,
(	71842	)	,
(	71876	)	,
(	71911	)	,
(	71945	)	,
(	71980	)	,
(	72014	)	,
(	72048	)	,
(	72083	)	,
(	72117	)	,
(	72152	)	,
(	72186	)	,
(	72221	)	,
(	72255	)	,
(	72290	)	,
(	72324	)	,
(	72359	)	,
(	72394	)	,
(	72428	)	,
(	72463	)	,
(	72497	)	,
(	72532	)	,
(	72567	)	,
(	72602	)	,
(	72636	)	,
(	72671	)	,
(	72706	)	,
(	72740	)	,
(	72775	)	,
(	72810	)	,
(	72845	)	,
(	72880	)	,
(	72915	)	,
(	72949	)	,
(	72984	)	,
(	73019	)	,
(	73054	)	,
(	73089	)	,
(	73124	)	,
(	73159	)	,
(	73194	)	,
(	73229	)	,
(	73264	)	,
(	73299	)	,
(	73334	)	,
(	73369	)	,
(	73404	)	,
(	73439	)	,
(	73474	)	,
(	73510	)	,
(	73545	)	,
(	73580	)	,
(	73615	)	,
(	73650	)	,
(	73685	)	,
(	73721	)	,
(	73756	)	,
(	73791	)	,
(	73826	)	,
(	73862	)	,
(	73897	)	,
(	73932	)	,
(	73968	)	,
(	74003	)	,
(	74039	)	,
(	74074	)	,
(	74109	)	,
(	74145	)	,
(	74180	)	,
(	74216	)	,
(	74251	)	,
(	74287	)	,
(	74322	)	,
(	74358	)	,
(	74393	)	,
(	74429	)	,
(	74464	)	,
(	74500	)	,
(	74536	)	,
(	74571	)	,
(	74607	)	,
(	74643	)	,
(	74678	)	,
(	74714	)	,
(	74750	)	,
(	74786	)	,
(	74821	)	,
(	74857	)	,
(	74893	)	,
(	74929	)	,
(	74964	)	,
(	75000	)	,
(	75036	)	,
(	75072	)	,
(	75108	)	,
(	75144	)	,
(	75180	)	,
(	75216	)	,
(	75252	)	,
(	75288	)	,
(	75324	)	,
(	75360	)	,
(	75396	)	,
(	75432	)	,
(	75468	)	,
(	75504	)	,
(	75540	)	,
(	75576	)	,
(	75612	)	,
(	75648	)	,
(	75685	)	,
(	75721	)	,
(	75757	)	,
(	75793	)	,
(	75829	)	,
(	75866	)	,
(	75902	)	,
(	75938	)	,
(	75975	)	,
(	76011	)	,
(	76047	)	,
(	76084	)	,
(	76120	)	,
(	76156	)	,
(	76193	)	,
(	76229	)	,
(	76266	)	,
(	76302	)	,
(	76339	)	,
(	76375	)	,
(	76412	)	,
(	76448	)	,
(	76485	)	,
(	76521	)	,
(	76558	)	,
(	76595	)	,
(	76631	)	,
(	76668	)	,
(	76704	)	,
(	76741	)	,
(	76778	)	,
(	76815	)	,
(	76851	)	,
(	76888	)	,
(	76925	)	,
(	76962	)	,
(	76998	)	,
(	77035	)	,
(	77072	)	,
(	77109	)	,
(	77146	)	,
(	77183	)	,
(	77220	)	,
(	77256	)	,
(	77293	)	,
(	77330	)	,
(	77367	)	,
(	77404	)	,
(	77441	)	,
(	77478	)	,
(	77515	)	,
(	77552	)	,
(	77590	)	,
(	77627	)	,
(	77664	)	,
(	77701	)	,
(	77738	)	,
(	77775	)	,
(	77812	)	,
(	77850	)	,
(	77887	)	,
(	77924	)	,
(	77961	)	,
(	77999	)	,
(	78036	)	,
(	78073	)	,
(	78111	)	,
(	78148	)	,
(	78185	)	,
(	78223	)	,
(	78260	)	,
(	78297	)	,
(	78335	)	,
(	78372	)	,
(	78410	)	,
(	78447	)	,
(	78485	)	,
(	78522	)	,
(	78560	)	,
(	78597	)	,
(	78635	)	,
(	78673	)	,
(	78710	)	,
(	78748	)	,
(	78786	)	,
(	78823	)	,
(	78861	)	,
(	78899	)	,
(	78936	)	,
(	78974	)	,
(	79012	)	,
(	79050	)	,
(	79087	)	,
(	79125	)	,
(	79163	)	,
(	79201	)	,
(	79239	)	,
(	79277	)	,
(	79315	)	,
(	79353	)	,
(	79390	)	,
(	79428	)	,
(	79466	)	,
(	79504	)	,
(	79542	)	,
(	79580	)	,
(	79618	)	,
(	79657	)	,
(	79695	)	,
(	79733	)	,
(	79771	)	,
(	79809	)	,
(	79847	)	,
(	79885	)	,
(	79924	)	,
(	79962	)	,
(	80000	)	,
(	80038	)	,
(	80077	)	,
(	80115	)	,
(	80153	)	,
(	80191	)	,
(	80230	)	,
(	80268	)	,
(	80307	)	,
(	80345	)	,
(	80383	)	,
(	80422	)	,
(	80460	)	,
(	80499	)	,
(	80537	)	,
(	80576	)	,
(	80614	)	,
(	80653	)	,
(	80691	)	,
(	80730	)	,
(	80769	)	,
(	80807	)	,
(	80846	)	,
(	80884	)	,
(	80923	)	,
(	80962	)	,
(	81001	)	,
(	81039	)	,
(	81078	)	,
(	81117	)	,
(	81156	)	,
(	81194	)	,
(	81233	)	,
(	81272	)	,
(	81311	)	,
(	81350	)	,
(	81389	)	,
(	81428	)	,
(	81466	)	,
(	81505	)	,
(	81544	)	,
(	81583	)	,
(	81622	)	,
(	81661	)	,
(	81700	)	,
(	81740	)	,
(	81779	)	,
(	81818	)	,
(	81857	)	,
(	81896	)	,
(	81935	)	,
(	81974	)	,
(	82014	)	,
(	82053	)	,
(	82092	)	,
(	82131	)	,
(	82171	)	,
(	82210	)	,
(	82249	)	,
(	82288	)	,
(	82328	)	,
(	82367	)	,
(	82407	)	,
(	82446	)	,
(	82485	)	,
(	82525	)	,
(	82564	)	,
(	82604	)	,
(	82643	)	,
(	82683	)	,
(	82722	)	,
(	82762	)	,
(	82801	)	,
(	82841	)	,
(	82881	)	,
(	82920	)	,
(	82960	)	,
(	83000	)	,
(	83039	)	,
(	83079	)	,
(	83119	)	,
(	83158	)	,
(	83198	)	,
(	83238	)	,
(	83278	)	,
(	83318	)	,
(	83357	)	,
(	83397	)	,
(	83437	)	,
(	83477	)	,
(	83517	)	,
(	83557	)	,
(	83597	)	,
(	83637	)	,
(	83677	)	,
(	83717	)	,
(	83757	)	,
(	83797	)	,
(	83837	)	,
(	83877	)	,
(	83917	)	,
(	83957	)	,
(	83997	)	,
(	84038	)	,
(	84078	)	,
(	84118	)	,
(	84158	)	,
(	84198	)	,
(	84239	)	,
(	84279	)	,
(	84319	)	,
(	84360	)	,
(	84400	)	,
(	84440	)	,
(	84481	)	,
(	84521	)	,
(	84561	)	,
(	84602	)	,
(	84642	)	,
(	84683	)	,
(	84723	)	,
(	84764	)	,
(	84804	)	,
(	84845	)	,
(	84885	)	,
(	84926	)	,
(	84967	)	,
(	85007	)	,
(	85048	)	,
(	85089	)	,
(	85129	)	,
(	85170	)	,
(	85211	)	,
(	85251	)	,
(	85292	)	,
(	85333	)	,
(	85374	)	,
(	85415	)	,
(	85455	)	,
(	85496	)	,
(	85537	)	,
(	85578	)	,
(	85619	)	,
(	85660	)	,
(	85701	)	,
(	85742	)	,
(	85783	)	,
(	85824	)	,
(	85865	)	,
(	85906	)	,
(	85947	)	,
(	85988	)	,
(	86029	)	,
(	86070	)	,
(	86112	)	,
(	86153	)	,
(	86194	)	,
(	86235	)	,
(	86276	)	,
(	86318	)	,
(	86359	)	,
(	86400	)	,
(	86442	)	,
(	86483	)	,
(	86524	)	,
(	86566	)	,
(	86607	)	,
(	86648	)	,
(	86690	)	,
(	86731	)	,
(	86773	)	,
(	86814	)	,
(	86856	)	,
(	86897	)	,
(	86939	)	,
(	86980	)	,
(	87022	)	,
(	87064	)	,
(	87105	)	,
(	87147	)	,
(	87189	)	,
(	87230	)	,
(	87272	)	,
(	87314	)	,
(	87355	)	,
(	87397	)	,
(	87439	)	,
(	87481	)	,
(	87523	)	,
(	87564	)	,
(	87606	)	,
(	87648	)	,
(	87690	)	,
(	87732	)	,
(	87774	)	,
(	87816	)	,
(	87858	)	,
(	87900	)	,
(	87942	)	,
(	87984	)	,
(	88026	)	,
(	88068	)	,
(	88110	)	,
(	88152	)	,
(	88195	)	,
(	88237	)	,
(	88279	)	,
(	88321	)	,
(	88363	)	,
(	88406	)	,
(	88448	)	,
(	88490	)	,
(	88532	)	,
(	88575	)	,
(	88617	)	,
(	88660	)	,
(	88702	)	,
(	88744	)	,
(	88787	)	,
(	88829	)	,
(	88872	)	,
(	88914	)	,
(	88957	)	,
(	88999	)	,
(	89042	)	,
(	89084	)	,
(	89127	)	,
(	89170	)	,
(	89212	)	,
(	89255	)	,
(	89298	)	,
(	89340	)	,
(	89383	)	,
(	89426	)	,
(	89468	)	,
(	89511	)	,
(	89554	)	,
(	89597	)	,
(	89640	)	,
(	89683	)	,
(	89725	)	,
(	89768	)	,
(	89811	)	,
(	89854	)	,
(	89897	)	,
(	89940	)	,
(	89983	)	,
(	90026	)	,
(	90069	)	,
(	90112	)	,
(	90155	)	,
(	90199	)	,
(	90242	)	,
(	90285	)	,
(	90328	)	,
(	90371	)	,
(	90414	)	,
(	90458	)	,
(	90501	)	,
(	90544	)	,
(	90587	)	,
(	90631	)	,
(	90674	)	,
(	90717	)	,
(	90761	)	,
(	90804	)	,
(	90848	)	,
(	90891	)	,
(	90934	)	,
(	90978	)	,
(	91021	)	,
(	91065	)	,
(	91109	)	,
(	91152	)	,
(	91196	)	,
(	91239	)	,
(	91283	)	,
(	91327	)	,
(	91370	)	,
(	91414	)	,
(	91458	)	,
(	91501	)	,
(	91545	)	,
(	91589	)	,
(	91633	)	,
(	91676	)	,
(	91720	)	,
(	91764	)	,
(	91808	)	,
(	91852	)	,
(	91896	)	,
(	91940	)	,
(	91984	)	,
(	92028	)	,
(	92072	)	,
(	92116	)	,
(	92160	)	,
(	92204	)	,
(	92248	)	,
(	92292	)	,
(	92336	)	,
(	92380	)	,
(	92425	)	,
(	92469	)	,
(	92513	)	,
(	92557	)	,
(	92601	)	,
(	92646	)	,
(	92690	)	,
(	92734	)	,
(	92779	)	,
(	92823	)	,
(	92867	)	,
(	92912	)	,
(	92956	)	,
(	93001	)	,
(	93045	)	,
(	93090	)	,
(	93134	)	,
(	93179	)	,
(	93223	)	,
(	93268	)	,
(	93312	)	,
(	93357	)	,
(	93402	)	,
(	93446	)	,
(	93491	)	,
(	93536	)	,
(	93580	)	,
(	93625	)	,
(	93670	)	,
(	93715	)	,
(	93760	)	,
(	93804	)	,
(	93849	)	,
(	93894	)	,
(	93939	)	,
(	93984	)	,
(	94029	)	,
(	94074	)	,
(	94119	)	,
(	94164	)	,
(	94209	)	,
(	94254	)	,
(	94299	)	,
(	94344	)	,
(	94389	)	,
(	94434	)	,
(	94479	)	,
(	94525	)	,
(	94570	)	,
(	94615	)	,
(	94660	)	,
(	94706	)	,
(	94751	)	,
(	94796	)	,
(	94841	)	,
(	94887	)	,
(	94932	)	,
(	94978	)	,
(	95023	)	,
(	95068	)	,
(	95114	)	,
(	95159	)	,
(	95205	)	,
(	95250	)	,
(	95296	)	,
(	95341	)	,
(	95387	)	,
(	95433	)	,
(	95478	)	,
(	95524	)	,
(	95570	)	,
(	95615	)	,
(	95661	)	,
(	95707	)	,
(	95753	)	,
(	95798	)	,
(	95844	)	,
(	95890	)	,
(	95936	)	,
(	95982	)	,
(	96028	)	,
(	96073	)	,
(	96119	)	,
(	96165	)	,
(	96211	)	,
(	96257	)	,
(	96303	)	,
(	96349	)	,
(	96395	)	,
(	96442	)	,
(	96488	)	,
(	96534	)	,
(	96580	)	,
(	96626	)	,
(	96672	)	,
(	96719	)	,
(	96765	)	,
(	96811	)	,
(	96857	)	,
(	96904	)	,
(	96950	)	,
(	96996	)	,
(	97043	)	,
(	97089	)	,
(	97136	)	,
(	97182	)	,
(	97229	)	,
(	97275	)	,
(	97322	)	,
(	97368	)	,
(	97415	)	,
(	97461	)	,
(	97508	)	,
(	97554	)	,
(	97601	)	,
(	97648	)	,
(	97694	)	,
(	97741	)	,
(	97788	)	,
(	97835	)	,
(	97881	)	,
(	97928	)	,
(	97975	)	,
(	98022	)	,
(	98069	)	,
(	98116	)	,
(	98163	)	,
(	98209	)	,
(	98256	)	,
(	98303	)	,
(	98350	)	,
(	98397	)	,
(	98444	)	,
(	98492	)	,
(	98539	)	,
(	98586	)	,
(	98633	)	,
(	98680	)	,
(	98727	)	,
(	98774	)	,
(	98822	)	,
(	98869	)	,
(	98916	)	,
(	98964	)	,
(	99011	)	,
(	99058	)	,
(	99106	)	,
(	99153	)	,
(	99200	)	,
(	99248	)	,
(	99295	)	,
(	99343	)	,
(	99390	)	,
(	99438	)	,
(	99485	)	,
(	99533	)	,
(	99580	)	,
(	99628	)	,
(	99676	)	,
(	99723	)	,
(	99771	)	,
(	99819	)	,
(	99866	)	,
(	99914	)	,
(	99962	)	,
(	100010	)	,
(	100058	)	,
(	100105	)	,
(	100153	)	,
(	100201	)	,
(	100249	)	,
(	100297	)	,
(	100345	)	,
(	100393	)	,
(	100441	)	,
(	100489	)	,
(	100537	)	,
(	100585	)	,
(	100633	)	,
(	100681	)	,
(	100729	)	,
(	100778	)	,
(	100826	)	,
(	100874	)	,
(	100922	)	,
(	100971	)	,
(	101019	)	,
(	101067	)	,
(	101115	)	,
(	101164	)	,
(	101212	)	,
(	101261	)	,
(	101309	)	,
(	101357	)	,
(	101406	)	,
(	101454	)	,
(	101503	)	,
(	101551	)	,
(	101600	)	,
(	101649	)	,
(	101697	)	,
(	101746	)	,
(	101794	)	,
(	101843	)	,
(	101892	)	,
(	101940	)	,
(	101989	)	,
(	102038	)	,
(	102087	)	,
(	102136	)	,
(	102184	)	,
(	102233	)	,
(	102282	)	,
(	102331	)	,
(	102380	)	,
(	102429	)	,
(	102478	)	,
(	102527	)	,
(	102576	)	,
(	102625	)	,
(	102674	)	,
(	102723	)	,
(	102772	)	,
(	102821	)	,
(	102871	)	,
(	102920	)	,
(	102969	)	,
(	103018	)	,
(	103067	)	,
(	103117	)	,
(	103166	)	,
(	103215	)	,
(	103265	)	,
(	103314	)	,
(	103364	)	,
(	103413	)	,
(	103462	)	,
(	103512	)	,
(	103561	)	,
(	103611	)	,
(	103660	)	,
(	103710	)	,
(	103760	)	,
(	103809	)	,
(	103859	)	,
(	103908	)	,
(	103958	)	,
(	104008	)	,
(	104058	)	,
(	104107	)	,
(	104157	)	,
(	104207	)	,
(	104257	)	,
(	104307	)	,
(	104356	)	,
(	104406	)	,
(	104456	)	,
(	104506	)	,
(	104556	)	,
(	104606	)	,
(	104656	)	,
(	104706	)	,
(	104756	)	,
(	104806	)	,
(	104857	)	,
(	104907	)	,
(	104957	)	,
(	105007	)	,
(	105057	)	,
(	105107	)	,
(	105158	)	,
(	105208	)	,
(	105258	)	,
(	105309	)	,
(	105359	)	,
(	105409	)	,
(	105460	)	,
(	105510	)	,
(	105561	)	,
(	105611	)	,
(	105662	)	,
(	105712	)	,
(	105763	)	,
(	105813	)	,
(	105864	)	,
(	105914	)	,
(	105965	)	,
(	106016	)	,
(	106066	)	,
(	106117	)	,
(	106168	)	,
(	106219	)	,
(	106269	)	,
(	106320	)	,
(	106371	)	,
(	106422	)	,
(	106473	)	,
(	106524	)	,
(	106575	)	,
(	106626	)	,
(	106677	)	,
(	106728	)	,
(	106779	)	,
(	106830	)	,
(	106881	)	,
(	106932	)	,
(	106983	)	,
(	107034	)	,
(	107085	)	,
(	107137	)	,
(	107188	)	,
(	107239	)	,
(	107290	)	,
(	107342	)	,
(	107393	)	,
(	107444	)	,
(	107496	)	,
(	107547	)	,
(	107599	)	,
(	107650	)	,
(	107701	)	,
(	107753	)	,
(	107804	)	,
(	107856	)	,
(	107908	)	,
(	107959	)	,
(	108011	)	,
(	108062	)	,
(	108114	)	,
(	108166	)	,
(	108218	)	,
(	108269	)	,
(	108321	)	,
(	108373	)	,
(	108425	)	,
(	108476	)	,
(	108528	)	,
(	108580	)	,
(	108632	)	,
(	108684	)	,
(	108736	)	,
(	108788	)	,
(	108840	)	,
(	108892	)	,
(	108944	)	,
(	108996	)	,
(	109048	)	,
(	109101	)	,
(	109153	)	,
(	109205	)	,
(	109257	)	,
(	109309	)	,
(	109362	)	,
(	109414	)	,
(	109466	)	,
(	109519	)	,
(	109571	)	,
(	109623	)	,
(	109676	)	,
(	109728	)	,
(	109781	)	,
(	109833	)	,
(	109886	)	,
(	109938	)	,
(	109991	)	,
(	110043	)	,
(	110096	)	,
(	110149	)	,
(	110201	)	,
(	110254	)	,
(	110307	)	,
(	110359	)	,
(	110412	)	,
(	110465	)	,
(	110518	)	,
(	110571	)	,
(	110624	)	,
(	110676	)	,
(	110729	)	,
(	110782	)	,
(	110835	)	,
(	110888	)	,
(	110941	)	,
(	110994	)	,
(	111047	)	,
(	111100	)	,
(	111154	)	,
(	111207	)	,
(	111260	)	,
(	111313	)	,
(	111366	)	,
(	111420	)	,
(	111473	)	,
(	111526	)	,
(	111579	)	,
(	111633	)	,
(	111686	)	,
(	111740	)	,
(	111793	)	,
(	111847	)	,
(	111900	)	,
(	111953	)	,
(	112007	)	,
(	112061	)	,
(	112114	)	,
(	112168	)	,
(	112221	)	,
(	112275	)	,
(	112329	)	,
(	112382	)	,
(	112436	)	,
(	112490	)	,
(	112544	)	,
(	112598	)	,
(	112651	)	,
(	112705	)	,
(	112759	)	,
(	112813	)	,
(	112867	)	,
(	112921	)	,
(	112975	)	,
(	113029	)	,
(	113083	)	,
(	113137	)	,
(	113191	)	,
(	113245	)	,
(	113299	)	,
(	113354	)	,
(	113408	)	,
(	113462	)	,
(	113516	)	,
(	113571	)	,
(	113625	)	,
(	113679	)	,
(	113734	)	,
(	113788	)	,
(	113842	)	,
(	113897	)	,
(	113951	)	,
(	114006	)	,
(	114060	)	,
(	114115	)	,
(	114169	)	,
(	114224	)	,
(	114279	)	,
(	114333	)	,
(	114388	)	,
(	114443	)	,
(	114497	)	,
(	114552	)	,
(	114607	)	,
(	114662	)	,
(	114716	)	,
(	114771	)	,
(	114826	)	,
(	114881	)	,
(	114936	)	,
(	114991	)	,
(	115046	)	,
(	115101	)	,
(	115156	)	,
(	115211	)	,
(	115266	)	,
(	115321	)	,
(	115376	)	,
(	115432	)	,
(	115487	)	,
(	115542	)	,
(	115597	)	,
(	115652	)	,
(	115708	)	,
(	115763	)	,
(	115818	)	,
(	115874	)	,
(	115929	)	,
(	115985	)	,
(	116040	)	,
(	116096	)	,
(	116151	)	,
(	116207	)	,
(	116262	)	,
(	116318	)	,
(	116373	)	,
(	116429	)	,
(	116485	)	,
(	116540	)	,
(	116596	)	,
(	116652	)	,
(	116708	)	,
(	116763	)	,
(	116819	)	,
(	116875	)	,
(	116931	)	,
(	116987	)	
	
);





begin
	
	determine_limit: process (clk, distance) is
	begin
		if rising_edge(clk) then
			if to_integer(unsigned(distance)) > 3300 then
				counter_limit <= to_unsigned(0, counter_limit'length);
			elsif to_integer(unsigned(distance)) < 0 then
				counter_limit <= to_unsigned(20000, counter_limit'length);
			else
				counter_limit <= to_unsigned(d2count(to_integer(unsigned(distance))),counter_limit'length);
			end if;
		end if;		
	end process;
	
	
	count: process (clk, reset) is
	begin		
		if rising_edge(clk) then
			if reset = '1' then
				counter <= to_unsigned(0, counter_limit'length);
			end if;
		
			counter <= counter + 1;
			
			if (counter > counter_limit) then
				counter <= to_unsigned(0, counter_limit'length);
			end if;
		end if;
	end process;
	

	produce_pwm : process(counter_limit, counter, reset)
   begin
		if reset = '1' or counter_limit = 0 then
			dac_out <= '0';
		else
			if (counter < (counter_limit / 2)) then  -- Potential issue unsigned(counter_limit)?
			  dac_out <= '0';
			else 
			  dac_out <= '1';
			end if;
		end if;
	end process;
				
end behavior;
