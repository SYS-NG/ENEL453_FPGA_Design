
-- In this example, we're going to map voltage to distance, using a linear 
-- approximation, according to the Sharp GP2Y0A41SK0F datasheet page 4, or 
-- Lab 3 handout page 5. 
-- 
-- The relevant points we will select are:
-- 2.750 V is  4.00 cm (or 2750 mV and  40.0 mm)
-- 0.400 V is 33.00 cm (or  400 mV and 330.0 mm)
-- 
-- Mapping to the scales in our system
-- 2750 (mV) should map to  400 (10^-4 m)
--  400 (mV) should map to 3300 (10^-4 m)
-- and developing a linear equation, we find:
--
-- Distance = -2900/2350 * Voltage + 3793.617
-- Note this code implements linear function, you must map to the 
-- NON-linear relationship in the datasheet. This code is only provided 
-- for reference to help get you started.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY voltage2distance IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;
		mux_bit_close  :  IN    STD_LOGIC;		
      voltage        :  IN    STD_LOGIC_VECTOR(12 DOWNTO 0);                           
      distance       :  OUT   STD_LOGIC_VECTOR(12 DOWNTO 0));
END voltage2distance;

ARCHITECTURE behavior OF voltage2distance IS

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.
-- See how to get the distance output at the bottom of this file,
-- after begin.

type array_1d is array (0 to 4095) of integer;
signal v_d_conversion : integer;

constant v2d_close: array_1d := (
(	-3	)	,
(	-3	)	,
(	-3	)	,
(	-3	)	,
(	-3	)	,
(	-2	)	,
(	-2	)	,
(	-2	)	,
(	-2	)	,
(	-2	)	,
(	-2	)	,
(	-2	)	,
(	-2	)	,
(	-2	)	,
(	-2	)	,
(	-1	)	,
(	-1	)	,
(	-1	)	,
(	-1	)	,
(	-1	)	,
(	-1	)	,
(	-1	)	,
(	-1	)	,
(	-1	)	,
(	-1	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	1	)	,
(	2	)	,
(	2	)	,
(	2	)	,
(	2	)	,
(	2	)	,
(	2	)	,
(	2	)	,
(	2	)	,
(	2	)	,
(	2	)	,
(	2	)	,
(	3	)	,
(	3	)	,
(	3	)	,
(	3	)	,
(	3	)	,
(	3	)	,
(	3	)	,
(	3	)	,
(	3	)	,
(	3	)	,
(	3	)	,
(	4	)	,
(	4	)	,
(	4	)	,
(	4	)	,
(	4	)	,
(	4	)	,
(	4	)	,
(	4	)	,
(	4	)	,
(	4	)	,
(	4	)	,
(	4	)	,
(	5	)	,
(	5	)	,
(	5	)	,
(	5	)	,
(	5	)	,
(	5	)	,
(	5	)	,
(	5	)	,
(	5	)	,
(	5	)	,
(	5	)	,
(	5	)	,
(	6	)	,
(	6	)	,
(	6	)	,
(	6	)	,
(	6	)	,
(	6	)	,
(	6	)	,
(	6	)	,
(	6	)	,
(	6	)	,
(	6	)	,
(	6	)	,
(	6	)	,
(	7	)	,
(	7	)	,
(	7	)	,
(	7	)	,
(	7	)	,
(	7	)	,
(	7	)	,
(	7	)	,
(	7	)	,
(	7	)	,
(	7	)	,
(	7	)	,
(	7	)	,
(	8	)	,
(	8	)	,
(	8	)	,
(	8	)	,
(	8	)	,
(	8	)	,
(	8	)	,
(	8	)	,
(	8	)	,
(	8	)	,
(	8	)	,
(	8	)	,
(	8	)	,
(	8	)	,
(	9	)	,
(	9	)	,
(	9	)	,
(	9	)	,
(	9	)	,
(	9	)	,
(	9	)	,
(	9	)	,
(	9	)	,
(	9	)	,
(	9	)	,
(	9	)	,
(	9	)	,
(	9	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	69	)	,
(	69	)	,
(	69	)	,
(	69	)	,
(	69	)	,
(	69	)	,
(	69	)	,
(	69	)	,
(	69	)	,
(	69	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	71	)	,
(	71	)	,
(	71	)	,
(	71	)	,
(	71	)	,
(	71	)	,
(	71	)	,
(	71	)	,
(	71	)	,
(	71	)	,
(	72	)	,
(	72	)	,
(	72	)	,
(	72	)	,
(	72	)	,
(	72	)	,
(	72	)	,
(	72	)	,
(	72	)	,
(	72	)	,
(	73	)	,
(	73	)	,
(	73	)	,
(	73	)	,
(	73	)	,
(	73	)	,
(	73	)	,
(	73	)	,
(	73	)	,
(	73	)	,
(	74	)	,
(	74	)	,
(	74	)	,
(	74	)	,
(	74	)	,
(	74	)	,
(	74	)	,
(	74	)	,
(	74	)	,
(	75	)	,
(	75	)	,
(	75	)	,
(	75	)	,
(	75	)	,
(	75	)	,
(	75	)	,
(	75	)	,
(	75	)	,
(	75	)	,
(	76	)	,
(	76	)	,
(	76	)	,
(	76	)	,
(	76	)	,
(	76	)	,
(	76	)	,
(	76	)	,
(	76	)	,
(	77	)	,
(	77	)	,
(	77	)	,
(	77	)	,
(	77	)	,
(	77	)	,
(	77	)	,
(	77	)	,
(	77	)	,
(	77	)	,
(	78	)	,
(	78	)	,
(	78	)	,
(	78	)	,
(	78	)	,
(	78	)	,
(	78	)	,
(	78	)	,
(	78	)	,
(	79	)	,
(	79	)	,
(	79	)	,
(	79	)	,
(	79	)	,
(	79	)	,
(	79	)	,
(	79	)	,
(	79	)	,
(	80	)	,
(	80	)	,
(	80	)	,
(	80	)	,
(	80	)	,
(	80	)	,
(	80	)	,
(	80	)	,
(	80	)	,
(	81	)	,
(	81	)	,
(	81	)	,
(	81	)	,
(	81	)	,
(	81	)	,
(	81	)	,
(	81	)	,
(	81	)	,
(	82	)	,
(	82	)	,
(	82	)	,
(	82	)	,
(	82	)	,
(	82	)	,
(	82	)	,
(	82	)	,
(	82	)	,
(	83	)	,
(	83	)	,
(	83	)	,
(	83	)	,
(	83	)	,
(	83	)	,
(	83	)	,
(	83	)	,
(	83	)	,
(	84	)	,
(	84	)	,
(	84	)	,
(	84	)	,
(	84	)	,
(	84	)	,
(	84	)	,
(	84	)	,
(	84	)	,
(	85	)	,
(	85	)	,
(	85	)	,
(	85	)	,
(	85	)	,
(	85	)	,
(	85	)	,
(	85	)	,
(	86	)	,
(	86	)	,
(	86	)	,
(	86	)	,
(	86	)	,
(	86	)	,
(	86	)	,
(	86	)	,
(	86	)	,
(	87	)	,
(	87	)	,
(	87	)	,
(	87	)	,
(	87	)	,
(	87	)	,
(	87	)	,
(	87	)	,
(	88	)	,
(	88	)	,
(	88	)	,
(	88	)	,
(	88	)	,
(	88	)	,
(	88	)	,
(	88	)	,
(	89	)	,
(	89	)	,
(	89	)	,
(	89	)	,
(	89	)	,
(	89	)	,
(	89	)	,
(	89	)	,
(	89	)	,
(	90	)	,
(	90	)	,
(	90	)	,
(	90	)	,
(	90	)	,
(	90	)	,
(	90	)	,
(	90	)	,
(	91	)	,
(	91	)	,
(	91	)	,
(	91	)	,
(	91	)	,
(	91	)	,
(	91	)	,
(	91	)	,
(	92	)	,
(	92	)	,
(	92	)	,
(	92	)	,
(	92	)	,
(	92	)	,
(	92	)	,
(	92	)	,
(	93	)	,
(	93	)	,
(	93	)	,
(	93	)	,
(	93	)	,
(	93	)	,
(	93	)	,
(	93	)	,
(	94	)	,
(	94	)	,
(	94	)	,
(	94	)	,
(	94	)	,
(	94	)	,
(	94	)	,
(	94	)	,
(	95	)	,
(	95	)	,
(	95	)	,
(	95	)	,
(	95	)	,
(	95	)	,
(	95	)	,
(	95	)	,
(	96	)	,
(	96	)	,
(	96	)	,
(	96	)	,
(	96	)	,
(	96	)	,
(	96	)	,
(	96	)	,
(	97	)	,
(	97	)	,
(	97	)	,
(	97	)	,
(	97	)	,
(	97	)	,
(	97	)	,
(	98	)	,
(	98	)	,
(	98	)	,
(	98	)	,
(	98	)	,
(	98	)	,
(	98	)	,
(	98	)	,
(	99	)	,
(	99	)	,
(	99	)	,
(	99	)	,
(	99	)	,
(	99	)	,
(	99	)	,
(	99	)	,
(	100	)	,
(	100	)	,
(	100	)	,
(	100	)	,
(	100	)	,
(	100	)	,
(	100	)	,
(	101	)	,
(	101	)	,
(	101	)	,
(	101	)	,
(	101	)	,
(	101	)	,
(	101	)	,
(	101	)	,
(	102	)	,
(	102	)	,
(	102	)	,
(	102	)	,
(	102	)	,
(	102	)	,
(	102	)	,
(	103	)	,
(	103	)	,
(	103	)	,
(	103	)	,
(	103	)	,
(	103	)	,
(	103	)	,
(	103	)	,
(	104	)	,
(	104	)	,
(	104	)	,
(	104	)	,
(	104	)	,
(	104	)	,
(	104	)	,
(	105	)	,
(	105	)	,
(	105	)	,
(	105	)	,
(	105	)	,
(	105	)	,
(	105	)	,
(	106	)	,
(	106	)	,
(	106	)	,
(	106	)	,
(	106	)	,
(	106	)	,
(	106	)	,
(	107	)	,
(	107	)	,
(	107	)	,
(	107	)	,
(	107	)	,
(	107	)	,
(	107	)	,
(	107	)	,
(	108	)	,
(	108	)	,
(	108	)	,
(	108	)	,
(	108	)	,
(	108	)	,
(	108	)	,
(	109	)	,
(	109	)	,
(	109	)	,
(	109	)	,
(	109	)	,
(	109	)	,
(	109	)	,
(	110	)	,
(	110	)	,
(	110	)	,
(	110	)	,
(	110	)	,
(	110	)	,
(	110	)	,
(	111	)	,
(	111	)	,
(	111	)	,
(	111	)	,
(	111	)	,
(	111	)	,
(	111	)	,
(	112	)	,
(	112	)	,
(	112	)	,
(	112	)	,
(	112	)	,
(	112	)	,
(	112	)	,
(	113	)	,
(	113	)	,
(	113	)	,
(	113	)	,
(	113	)	,
(	113	)	,
(	113	)	,
(	114	)	,
(	114	)	,
(	114	)	,
(	114	)	,
(	114	)	,
(	114	)	,
(	114	)	,
(	115	)	,
(	115	)	,
(	115	)	,
(	115	)	,
(	115	)	,
(	115	)	,
(	115	)	,
(	116	)	,
(	116	)	,
(	116	)	,
(	116	)	,
(	116	)	,
(	116	)	,
(	117	)	,
(	117	)	,
(	117	)	,
(	117	)	,
(	117	)	,
(	117	)	,
(	117	)	,
(	118	)	,
(	118	)	,
(	118	)	,
(	118	)	,
(	118	)	,
(	118	)	,
(	118	)	,
(	119	)	,
(	119	)	,
(	119	)	,
(	119	)	,
(	119	)	,
(	119	)	,
(	119	)	,
(	120	)	,
(	120	)	,
(	120	)	,
(	120	)	,
(	120	)	,
(	120	)	,
(	121	)	,
(	121	)	,
(	121	)	,
(	121	)	,
(	121	)	,
(	121	)	,
(	121	)	,
(	122	)	,
(	122	)	,
(	122	)	,
(	122	)	,
(	122	)	,
(	122	)	,
(	123	)	,
(	123	)	,
(	123	)	,
(	123	)	,
(	123	)	,
(	123	)	,
(	123	)	,
(	124	)	,
(	124	)	,
(	124	)	,
(	124	)	,
(	124	)	,
(	124	)	,
(	124	)	,
(	125	)	,
(	125	)	,
(	125	)	,
(	125	)	,
(	125	)	,
(	125	)	,
(	126	)	,
(	126	)	,
(	126	)	,
(	126	)	,
(	126	)	,
(	126	)	,
(	127	)	,
(	127	)	,
(	127	)	,
(	127	)	,
(	127	)	,
(	127	)	,
(	127	)	,
(	128	)	,
(	128	)	,
(	128	)	,
(	128	)	,
(	128	)	,
(	128	)	,
(	129	)	,
(	129	)	,
(	129	)	,
(	129	)	,
(	129	)	,
(	129	)	,
(	129	)	,
(	130	)	,
(	130	)	,
(	130	)	,
(	130	)	,
(	130	)	,
(	130	)	,
(	131	)	,
(	131	)	,
(	131	)	,
(	131	)	,
(	131	)	,
(	131	)	,
(	132	)	,
(	132	)	,
(	132	)	,
(	132	)	,
(	132	)	,
(	132	)	,
(	132	)	,
(	133	)	,
(	133	)	,
(	133	)	,
(	133	)	,
(	133	)	,
(	133	)	,
(	134	)	,
(	134	)	,
(	134	)	,
(	134	)	,
(	134	)	,
(	134	)	,
(	135	)	,
(	135	)	,
(	135	)	,
(	135	)	,
(	135	)	,
(	135	)	,
(	136	)	,
(	136	)	,
(	136	)	,
(	136	)	,
(	136	)	,
(	136	)	,
(	136	)	,
(	137	)	,
(	137	)	,
(	137	)	,
(	137	)	,
(	137	)	,
(	137	)	,
(	138	)	,
(	138	)	,
(	138	)	,
(	138	)	,
(	138	)	,
(	138	)	,
(	139	)	,
(	139	)	,
(	139	)	,
(	139	)	,
(	139	)	,
(	139	)	,
(	140	)	,
(	140	)	,
(	140	)	,
(	140	)	,
(	140	)	,
(	140	)	,
(	141	)	,
(	141	)	,
(	141	)	,
(	141	)	,
(	141	)	,
(	141	)	,
(	142	)	,
(	142	)	,
(	142	)	,
(	142	)	,
(	142	)	,
(	142	)	,
(	143	)	,
(	143	)	,
(	143	)	,
(	143	)	,
(	143	)	,
(	143	)	,
(	144	)	,
(	144	)	,
(	144	)	,
(	144	)	,
(	144	)	,
(	144	)	,
(	145	)	,
(	145	)	,
(	145	)	,
(	145	)	,
(	145	)	,
(	145	)	,
(	146	)	,
(	146	)	,
(	146	)	,
(	146	)	,
(	146	)	,
(	146	)	,
(	147	)	,
(	147	)	,
(	147	)	,
(	147	)	,
(	147	)	,
(	147	)	,
(	148	)	,
(	148	)	,
(	148	)	,
(	148	)	,
(	148	)	,
(	148	)	,
(	149	)	,
(	149	)	,
(	149	)	,
(	149	)	,
(	149	)	,
(	149	)	,
(	150	)	,
(	150	)	,
(	150	)	,
(	150	)	,
(	150	)	,
(	150	)	,
(	151	)	,
(	151	)	,
(	151	)	,
(	151	)	,
(	151	)	,
(	151	)	,
(	152	)	,
(	152	)	,
(	152	)	,
(	152	)	,
(	152	)	,
(	153	)	,
(	153	)	,
(	153	)	,
(	153	)	,
(	153	)	,
(	153	)	,
(	154	)	,
(	154	)	,
(	154	)	,
(	154	)	,
(	154	)	,
(	154	)	,
(	155	)	,
(	155	)	,
(	155	)	,
(	155	)	,
(	155	)	,
(	155	)	,
(	156	)	,
(	156	)	,
(	156	)	,
(	156	)	,
(	156	)	,
(	156	)	,
(	157	)	,
(	157	)	,
(	157	)	,
(	157	)	,
(	157	)	,
(	158	)	,
(	158	)	,
(	158	)	,
(	158	)	,
(	158	)	,
(	158	)	,
(	159	)	,
(	159	)	,
(	159	)	,
(	159	)	,
(	159	)	,
(	159	)	,
(	160	)	,
(	160	)	,
(	160	)	,
(	160	)	,
(	160	)	,
(	160	)	,
(	161	)	,
(	161	)	,
(	161	)	,
(	161	)	,
(	161	)	,
(	162	)	,
(	162	)	,
(	162	)	,
(	162	)	,
(	162	)	,
(	162	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	164	)	,
(	164	)	,
(	164	)	,
(	164	)	,
(	164	)	,
(	165	)	,
(	165	)	,
(	165	)	,
(	165	)	,
(	165	)	,
(	165	)	,
(	166	)	,
(	166	)	,
(	166	)	,
(	166	)	,
(	166	)	,
(	166	)	,
(	167	)	,
(	167	)	,
(	167	)	,
(	167	)	,
(	167	)	,
(	168	)	,
(	168	)	,
(	168	)	,
(	168	)	,
(	168	)	,
(	168	)	,
(	169	)	,
(	169	)	,
(	169	)	,
(	169	)	,
(	169	)	,
(	170	)	,
(	170	)	,
(	170	)	,
(	170	)	,
(	170	)	,
(	170	)	,
(	171	)	,
(	171	)	,
(	171	)	,
(	171	)	,
(	171	)	,
(	172	)	,
(	172	)	,
(	172	)	,
(	172	)	,
(	172	)	,
(	172	)	,
(	173	)	,
(	173	)	,
(	173	)	,
(	173	)	,
(	173	)	,
(	174	)	,
(	174	)	,
(	174	)	,
(	174	)	,
(	174	)	,
(	174	)	,
(	175	)	,
(	175	)	,
(	175	)	,
(	175	)	,
(	175	)	,
(	175	)	,
(	176	)	,
(	176	)	,
(	176	)	,
(	176	)	,
(	176	)	,
(	177	)	,
(	177	)	,
(	177	)	,
(	177	)	,
(	177	)	,
(	178	)	,
(	178	)	,
(	178	)	,
(	178	)	,
(	178	)	,
(	178	)	,
(	179	)	,
(	179	)	,
(	179	)	,
(	179	)	,
(	179	)	,
(	180	)	,
(	180	)	,
(	180	)	,
(	180	)	,
(	180	)	,
(	180	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	181	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	182	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	183	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	184	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	185	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	186	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	187	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	188	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	189	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	190	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	191	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	192	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	193	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	194	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	195	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	196	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	197	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	198	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	199	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	200	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	201	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	202	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	203	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	204	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	205	)	,
(	206	)	,
(	206	)	,
(	206	)	,
(	206	)	,
(	206	)	,
(	206	)	,
(	207	)	,
(	207	)	,
(	207	)	,
(	207	)	,
(	207	)	,
(	208	)	,
(	208	)	,
(	208	)	,
(	208	)	,
(	208	)	,
(	209	)	,
(	209	)	,
(	209	)	,
(	209	)	,
(	209	)	,
(	210	)	,
(	210	)	,
(	210	)	,
(	210	)	,
(	210	)	,
(	210	)	,
(	211	)	,
(	211	)	,
(	211	)	,
(	211	)	,
(	211	)	,
(	212	)	,
(	212	)	,
(	212	)	,
(	212	)	,
(	212	)	,
(	213	)	,
(	213	)	,
(	213	)	,
(	213	)	,
(	213	)	,
(	214	)	,
(	214	)	,
(	214	)	,
(	214	)	,
(	214	)	,
(	214	)	,
(	215	)	,
(	215	)	,
(	215	)	,
(	215	)	,
(	215	)	,
(	216	)	,
(	216	)	,
(	216	)	,
(	216	)	,
(	216	)	,
(	217	)	,
(	217	)	,
(	217	)	,
(	217	)	,
(	217	)	,
(	218	)	,
(	218	)	,
(	218	)	,
(	218	)	,
(	218	)	,
(	218	)	,
(	219	)	,
(	219	)	,
(	219	)	,
(	219	)	,
(	219	)	,
(	220	)	,
(	220	)	,
(	220	)	,
(	220	)	,
(	220	)	,
(	221	)	,
(	221	)	,
(	221	)	,
(	221	)	,
(	221	)	,
(	222	)	,
(	222	)	,
(	222	)	,
(	222	)	,
(	222	)	,
(	223	)	,
(	223	)	,
(	223	)	,
(	223	)	,
(	223	)	,
(	223	)	,
(	224	)	,
(	224	)	,
(	224	)	,
(	224	)	,
(	224	)	,
(	225	)	,
(	225	)	,
(	225	)	,
(	225	)	,
(	225	)	,
(	226	)	,
(	226	)	,
(	226	)	,
(	226	)	,
(	226	)	,
(	227	)	,
(	227	)	,
(	227	)	,
(	227	)	,
(	227	)	,
(	228	)	,
(	228	)	,
(	228	)	,
(	228	)	,
(	228	)	,
(	228	)	,
(	229	)	,
(	229	)	,
(	229	)	,
(	229	)	,
(	229	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	230	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	231	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	232	)	,
(	233	)	,
(	233	)	,
(	233	)	,
(	233	)	,
(	233	)	,
(	234	)	,
(	234	)	,
(	234	)	,
(	234	)	,
(	234	)	,
(	235	)	,
(	235	)	,
(	235	)	,
(	235	)	,
(	235	)	,
(	236	)	,
(	236	)	,
(	236	)	,
(	236	)	,
(	236	)	,
(	237	)	,
(	237	)	,
(	237	)	,
(	237	)	,
(	237	)	,
(	237	)	,
(	238	)	,
(	238	)	,
(	238	)	,
(	238	)	,
(	238	)	,
(	239	)	,
(	239	)	,
(	239	)	,
(	239	)	,
(	239	)	,
(	240	)	,
(	240	)	,
(	240	)	,
(	240	)	,
(	240	)	,
(	241	)	,
(	241	)	,
(	241	)	,
(	241	)	,
(	241	)	,
(	242	)	,
(	242	)	,
(	242	)	,
(	242	)	,
(	242	)	,
(	242	)	,
(	243	)	,
(	243	)	,
(	243	)	,
(	243	)	,
(	243	)	,
(	244	)	,
(	244	)	,
(	244	)	,
(	244	)	,
(	244	)	,
(	245	)	,
(	245	)	,
(	245	)	,
(	245	)	,
(	245	)	,
(	246	)	,
(	246	)	,
(	246	)	,
(	246	)	,
(	246	)	,
(	246	)	,
(	247	)	,
(	247	)	,
(	247	)	,
(	247	)	,
(	247	)	,
(	248	)	,
(	248	)	,
(	248	)	,
(	248	)	,
(	248	)	,
(	249	)	,
(	249	)	,
(	249	)	,
(	249	)	,
(	249	)	,
(	250	)	,
(	250	)	,
(	250	)	,
(	250	)	,
(	250	)	,
(	250	)	,
(	251	)	,
(	251	)	,
(	251	)	,
(	251	)	,
(	251	)	,
(	252	)	,
(	252	)	,
(	252	)	,
(	252	)	,
(	252	)	,
(	253	)	,
(	253	)	,
(	253	)	,
(	253	)	,
(	253	)	,
(	253	)	,
(	254	)	,
(	254	)	,
(	254	)	,
(	254	)	,
(	254	)	,
(	255	)	,
(	255	)	,
(	255	)	,
(	255	)	,
(	255	)	,
(	256	)	,
(	256	)	,
(	256	)	,
(	256	)	,
(	256	)	,
(	257	)	,
(	257	)	,
(	257	)	,
(	257	)	,
(	257	)	,
(	257	)	,
(	258	)	,
(	258	)	,
(	258	)	,
(	258	)	,
(	258	)	,
(	259	)	,
(	259	)	,
(	259	)	,
(	259	)	,
(	259	)	,
(	260	)	,
(	260	)	,
(	260	)	,
(	260	)	,
(	260	)	,
(	260	)	,
(	261	)	,
(	261	)	,
(	261	)	,
(	261	)	,
(	261	)	,
(	262	)	,
(	262	)	,
(	262	)	,
(	262	)	,
(	262	)	,
(	263	)	,
(	263	)	,
(	263	)	,
(	263	)	,
(	263	)	,
(	263	)	,
(	264	)	,
(	264	)	,
(	264	)	,
(	264	)	,
(	264	)	,
(	265	)	,
(	265	)	,
(	265	)	,
(	265	)	,
(	265	)	,
(	266	)	,
(	266	)	,
(	266	)	,
(	266	)	,
(	266	)	,
(	266	)	,
(	267	)	,
(	267	)	,
(	267	)	,
(	267	)	,
(	267	)	,
(	268	)	,
(	268	)	,
(	268	)	,
(	268	)	,
(	268	)	,
(	268	)	,
(	269	)	,
(	269	)	,
(	269	)	,
(	269	)	,
(	269	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	273	)	,
(	273	)	,
(	273	)	,
(	273	)	,
(	273	)	,
(	273	)	,
(	274	)	,
(	274	)	,
(	274	)	,
(	274	)	,
(	274	)	,
(	275	)	,
(	275	)	,
(	275	)	,
(	275	)	,
(	275	)	,
(	275	)	,
(	276	)	,
(	276	)	,
(	276	)	,
(	276	)	,
(	276	)	,
(	277	)	,
(	277	)	,
(	277	)	,
(	277	)	,
(	277	)	,
(	277	)	,
(	278	)	,
(	278	)	,
(	278	)	,
(	278	)	,
(	278	)	,
(	279	)	,
(	279	)	,
(	279	)	,
(	279	)	,
(	279	)	,
(	279	)	,
(	280	)	,
(	280	)	,
(	280	)	,
(	280	)	,
(	280	)	,
(	281	)	,
(	281	)	,
(	281	)	,
(	281	)	,
(	281	)	,
(	281	)	,
(	282	)	,
(	282	)	,
(	282	)	,
(	282	)	,
(	282	)	,
(	283	)	,
(	283	)	,
(	283	)	,
(	283	)	,
(	283	)	,
(	283	)	,
(	284	)	,
(	284	)	,
(	284	)	,
(	284	)	,
(	284	)	,
(	284	)	,
(	285	)	,
(	285	)	,
(	285	)	,
(	285	)	,
(	285	)	,
(	286	)	,
(	286	)	,
(	286	)	,
(	286	)	,
(	286	)	,
(	286	)	,
(	287	)	,
(	287	)	,
(	287	)	,
(	287	)	,
(	287	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	292	)	,
(	292	)	,
(	292	)	,
(	292	)	,
(	292	)	,
(	292	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	294	)	,
(	295	)	,
(	295	)	,
(	295	)	,
(	295	)	,
(	295	)	,
(	295	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	297	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	299	)	,
(	299	)	,
(	299	)	,
(	299	)	,
(	299	)	,
(	299	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	300	)	,
(	301	)	,
(	301	)	,
(	301	)	,
(	301	)	,
(	301	)	,
(	301	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	302	)	,
(	303	)	,
(	303	)	,
(	303	)	,
(	303	)	,
(	303	)	,
(	303	)	,
(	304	)	,
(	304	)	,
(	304	)	,
(	304	)	,
(	304	)	,
(	304	)	,
(	305	)	,
(	305	)	,
(	305	)	,
(	305	)	,
(	305	)	,
(	305	)	,
(	306	)	,
(	306	)	,
(	306	)	,
(	306	)	,
(	306	)	,
(	306	)	,
(	307	)	,
(	307	)	,
(	307	)	,
(	307	)	,
(	307	)	,
(	307	)	,
(	307	)	,
(	308	)	,
(	308	)	,
(	308	)	,
(	308	)	,
(	308	)	,
(	308	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	316	)	,
(	316	)	,
(	316	)	,
(	316	)	,
(	316	)	,
(	316	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	318	)	,
(	318	)	,
(	318	)	,
(	318	)	,
(	318	)	,
(	318	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	361	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	360	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	359	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	358	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	357	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	356	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	355	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	354	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	353	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	352	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	351	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	350	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	349	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	348	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	347	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	346	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	345	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	344	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	343	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	342	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	341	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	340	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	339	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	338	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	337	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	336	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	335	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	334	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	333	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	332	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	331	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	330	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	329	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	328	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	327	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	326	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	325	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	324	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	323	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	322	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	321	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	320	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	319	)	,
(	318	)	,
(	318	)	,
(	318	)	,
(	318	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	317	)	,
(	316	)	,
(	316	)	,
(	316	)	,
(	316	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	315	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	314	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	313	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	312	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	311	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	310	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	309	)	,
(	308	)	,
(	308	)	,
(	308	)	
);

constant v2d_LUT : array_1d := (

(	8343	)	,
(	8324	)	,
(	8305	)	,
(	8286	)	,
(	8267	)	,
(	8248	)	,
(	8229	)	,
(	8210	)	,
(	8191	)	,
(	8172	)	,
(	8154	)	,
(	8135	)	,
(	8116	)	,
(	8098	)	,
(	8079	)	,
(	8060	)	,
(	8042	)	,
(	8023	)	,
(	8005	)	,
(	7987	)	,
(	7968	)	,
(	7950	)	,
(	7932	)	,
(	7913	)	,
(	7895	)	,
(	7877	)	,
(	7859	)	,
(	7841	)	,
(	7823	)	,
(	7805	)	,
(	7787	)	,
(	7769	)	,
(	7751	)	,
(	7733	)	,
(	7715	)	,
(	7697	)	,
(	7680	)	,
(	7662	)	,
(	7644	)	,
(	7627	)	,
(	7609	)	,
(	7592	)	,
(	7574	)	,
(	7557	)	,
(	7539	)	,
(	7522	)	,
(	7504	)	,
(	7487	)	,
(	7470	)	,
(	7453	)	,
(	7435	)	,
(	7418	)	,
(	7401	)	,
(	7384	)	,
(	7367	)	,
(	7350	)	,
(	7333	)	,
(	7316	)	,
(	7299	)	,
(	7282	)	,
(	7266	)	,
(	7249	)	,
(	7232	)	,
(	7215	)	,
(	7199	)	,
(	7182	)	,
(	7165	)	,
(	7149	)	,
(	7132	)	,
(	7116	)	,
(	7099	)	,
(	7083	)	,
(	7067	)	,
(	7050	)	,
(	7034	)	,
(	7018	)	,
(	7001	)	,
(	6985	)	,
(	6969	)	,
(	6953	)	,
(	6937	)	,
(	6921	)	,
(	6905	)	,
(	6889	)	,
(	6873	)	,
(	6857	)	,
(	6841	)	,
(	6825	)	,
(	6810	)	,
(	6794	)	,
(	6778	)	,
(	6762	)	,
(	6747	)	,
(	6731	)	,
(	6716	)	,
(	6700	)	,
(	6684	)	,
(	6669	)	,
(	6654	)	,
(	6638	)	,
(	6623	)	,
(	6607	)	,
(	6592	)	,
(	6577	)	,
(	6562	)	,
(	6546	)	,
(	6531	)	,
(	6516	)	,
(	6501	)	,
(	6486	)	,
(	6471	)	,
(	6456	)	,
(	6441	)	,
(	6426	)	,
(	6411	)	,
(	6396	)	,
(	6382	)	,
(	6367	)	,
(	6352	)	,
(	6337	)	,
(	6323	)	,
(	6308	)	,
(	6293	)	,
(	6279	)	,
(	6264	)	,
(	6250	)	,
(	6235	)	,
(	6221	)	,
(	6206	)	,
(	6192	)	,
(	6178	)	,
(	6163	)	,
(	6149	)	,
(	6135	)	,
(	6121	)	,
(	6106	)	,
(	6092	)	,
(	6078	)	,
(	6064	)	,
(	6050	)	,
(	6036	)	,
(	6022	)	,
(	6008	)	,
(	5994	)	,
(	5980	)	,
(	5966	)	,
(	5952	)	,
(	5939	)	,
(	5925	)	,
(	5911	)	,
(	5897	)	,
(	5884	)	,
(	5870	)	,
(	5857	)	,
(	5843	)	,
(	5829	)	,
(	5816	)	,
(	5802	)	,
(	5789	)	,
(	5776	)	,
(	5762	)	,
(	5749	)	,
(	5736	)	,
(	5722	)	,
(	5709	)	,
(	5696	)	,
(	5683	)	,
(	5669	)	,
(	5656	)	,
(	5643	)	,
(	5630	)	,
(	5617	)	,
(	5604	)	,
(	5591	)	,
(	5578	)	,
(	5565	)	,
(	5552	)	,
(	5540	)	,
(	5527	)	,
(	5514	)	,
(	5501	)	,
(	5488	)	,
(	5476	)	,
(	5463	)	,
(	5450	)	,
(	5438	)	,
(	5425	)	,
(	5413	)	,
(	5400	)	,
(	5388	)	,
(	5375	)	,
(	5363	)	,
(	5350	)	,
(	5338	)	,
(	5326	)	,
(	5313	)	,
(	5301	)	,
(	5289	)	,
(	5277	)	,
(	5264	)	,
(	5252	)	,
(	5240	)	,
(	5228	)	,
(	5216	)	,
(	5204	)	,
(	5192	)	,
(	5180	)	,
(	5168	)	,
(	5156	)	,
(	5144	)	,
(	5132	)	,
(	5120	)	,
(	5108	)	,
(	5097	)	,
(	5085	)	,
(	5073	)	,
(	5061	)	,
(	5050	)	,
(	5038	)	,
(	5026	)	,
(	5015	)	,
(	5003	)	,
(	4992	)	,
(	4980	)	,
(	4969	)	,
(	4957	)	,
(	4946	)	,
(	4934	)	,
(	4923	)	,
(	4912	)	,
(	4900	)	,
(	4889	)	,
(	4878	)	,
(	4867	)	,
(	4855	)	,
(	4844	)	,
(	4833	)	,
(	4822	)	,
(	4811	)	,
(	4800	)	,
(	4789	)	,
(	4778	)	,
(	4767	)	,
(	4756	)	,
(	4745	)	,
(	4734	)	,
(	4723	)	,
(	4712	)	,
(	4701	)	,
(	4691	)	,
(	4680	)	,
(	4669	)	,
(	4658	)	,
(	4648	)	,
(	4637	)	,
(	4626	)	,
(	4616	)	,
(	4605	)	,
(	4595	)	,
(	4584	)	,
(	4574	)	,
(	4563	)	,
(	4553	)	,
(	4542	)	,
(	4532	)	,
(	4521	)	,
(	4511	)	,
(	4501	)	,
(	4490	)	,
(	4480	)	,
(	4470	)	,
(	4460	)	,
(	4449	)	,
(	4439	)	,
(	4429	)	,
(	4419	)	,
(	4409	)	,
(	4399	)	,
(	4389	)	,
(	4379	)	,
(	4369	)	,
(	4359	)	,
(	4349	)	,
(	4339	)	,
(	4329	)	,
(	4319	)	,
(	4309	)	,
(	4299	)	,
(	4290	)	,
(	4280	)	,
(	4270	)	,
(	4260	)	,
(	4251	)	,
(	4241	)	,
(	4231	)	,
(	4222	)	,
(	4212	)	,
(	4202	)	,
(	4193	)	,
(	4183	)	,
(	4174	)	,
(	4164	)	,
(	4155	)	,
(	4145	)	,
(	4136	)	,
(	4127	)	,
(	4117	)	,
(	4108	)	,
(	4099	)	,
(	4089	)	,
(	4080	)	,
(	4071	)	,
(	4062	)	,
(	4052	)	,
(	4043	)	,
(	4034	)	,
(	4025	)	,
(	4016	)	,
(	4007	)	,
(	3998	)	,
(	3989	)	,
(	3980	)	,
(	3971	)	,
(	3962	)	,
(	3953	)	,
(	3944	)	,
(	3935	)	,
(	3926	)	,
(	3917	)	,
(	3908	)	,
(	3900	)	,
(	3891	)	,
(	3882	)	,
(	3873	)	,
(	3865	)	,
(	3856	)	,
(	3847	)	,
(	3839	)	,
(	3830	)	,
(	3821	)	,
(	3813	)	,
(	3804	)	,
(	3796	)	,
(	3787	)	,
(	3779	)	,
(	3770	)	,
(	3762	)	,
(	3753	)	,
(	3745	)	,
(	3736	)	,
(	3728	)	,
(	3720	)	,
(	3711	)	,
(	3703	)	,
(	3695	)	,
(	3687	)	,
(	3678	)	,
(	3670	)	,
(	3662	)	,
(	3654	)	,
(	3646	)	,
(	3638	)	,
(	3629	)	,
(	3621	)	,
(	3613	)	,
(	3605	)	,
(	3597	)	,
(	3589	)	,
(	3581	)	,
(	3573	)	,
(	3565	)	,
(	3557	)	,
(	3550	)	,
(	3542	)	,
(	3534	)	,
(	3526	)	,
(	3518	)	,
(	3510	)	,
(	3503	)	,
(	3495	)	,
(	3487	)	,
(	3479	)	,
(	3472	)	,
(	3464	)	,
(	3456	)	,
(	3449	)	,
(	3441	)	,
(	3434	)	,
(	3426	)	,
(	3419	)	,
(	3411	)	,
(	3404	)	,
(	3396	)	,
(	3389	)	,
(	3381	)	,
(	3374	)	,
(	3366	)	,
(	3359	)	,
(	3352	)	,
(	3344	)	,
(	3337	)	,
(	3330	)	,
(	3322	)	,
(	3315	)	,
(	3308	)	,
(	3300	)	,
(	3293	)	,
(	3286	)	,
(	3279	)	,
(	3272	)	,
(	3265	)	,
(	3258	)	,
(	3250	)	,
(	3243	)	,
(	3236	)	,
(	3229	)	,
(	3222	)	,
(	3215	)	,
(	3208	)	,
(	3201	)	,
(	3194	)	,
(	3187	)	,
(	3181	)	,
(	3174	)	,
(	3167	)	,
(	3160	)	,
(	3153	)	,
(	3146	)	,
(	3139	)	,
(	3133	)	,
(	3126	)	,
(	3119	)	,
(	3112	)	,
(	3106	)	,
(	3099	)	,
(	3092	)	,
(	3086	)	,
(	3079	)	,
(	3073	)	,
(	3066	)	,
(	3059	)	,
(	3053	)	,
(	3046	)	,
(	3040	)	,
(	3033	)	,
(	3027	)	,
(	3020	)	,
(	3014	)	,
(	3007	)	,
(	3001	)	,
(	2995	)	,
(	2988	)	,
(	2982	)	,
(	2975	)	,
(	2969	)	,
(	2963	)	,
(	2957	)	,
(	2950	)	,
(	2944	)	,
(	2938	)	,
(	2932	)	,
(	2925	)	,
(	2919	)	,
(	2913	)	,
(	2907	)	,
(	2901	)	,
(	2895	)	,
(	2888	)	,
(	2882	)	,
(	2876	)	,
(	2870	)	,
(	2864	)	,
(	2858	)	,
(	2852	)	,
(	2846	)	,
(	2840	)	,
(	2834	)	,
(	2828	)	,
(	2822	)	,
(	2816	)	,
(	2811	)	,
(	2805	)	,
(	2799	)	,
(	2793	)	,
(	2787	)	,
(	2781	)	,
(	2776	)	,
(	2770	)	,
(	2764	)	,
(	2758	)	,
(	2753	)	,
(	2747	)	,
(	2741	)	,
(	2736	)	,
(	2730	)	,
(	2724	)	,
(	2719	)	,
(	2713	)	,
(	2707	)	,
(	2702	)	,
(	2696	)	,
(	2691	)	,
(	2685	)	,
(	2680	)	,
(	2674	)	,
(	2669	)	,
(	2663	)	,
(	2658	)	,
(	2652	)	,
(	2647	)	,
(	2641	)	,
(	2636	)	,
(	2631	)	,
(	2625	)	,
(	2620	)	,
(	2615	)	,
(	2609	)	,
(	2604	)	,
(	2599	)	,
(	2593	)	,
(	2588	)	,
(	2583	)	,
(	2578	)	,
(	2572	)	,
(	2567	)	,
(	2562	)	,
(	2557	)	,
(	2552	)	,
(	2547	)	,
(	2541	)	,
(	2536	)	,
(	2531	)	,
(	2526	)	,
(	2521	)	,
(	2516	)	,
(	2511	)	,
(	2506	)	,
(	2501	)	,
(	2496	)	,
(	2491	)	,
(	2486	)	,
(	2481	)	,
(	2476	)	,
(	2471	)	,
(	2466	)	,
(	2461	)	,
(	2457	)	,
(	2452	)	,
(	2447	)	,
(	2442	)	,
(	2437	)	,
(	2432	)	,
(	2428	)	,
(	2423	)	,
(	2418	)	,
(	2413	)	,
(	2408	)	,
(	2404	)	,
(	2399	)	,
(	2394	)	,
(	2390	)	,
(	2385	)	,
(	2380	)	,
(	2376	)	,
(	2371	)	,
(	2366	)	,
(	2362	)	,
(	2357	)	,
(	2353	)	,
(	2348	)	,
(	2344	)	,
(	2339	)	,
(	2334	)	,
(	2330	)	,
(	2325	)	,
(	2321	)	,
(	2316	)	,
(	2312	)	,
(	2308	)	,
(	2303	)	,
(	2299	)	,
(	2294	)	,
(	2290	)	,
(	2286	)	,
(	2281	)	,
(	2277	)	,
(	2272	)	,
(	2268	)	,
(	2264	)	,
(	2259	)	,
(	2255	)	,
(	2251	)	,
(	2247	)	,
(	2242	)	,
(	2238	)	,
(	2234	)	,
(	2230	)	,
(	2225	)	,
(	2221	)	,
(	2217	)	,
(	2213	)	,
(	2209	)	,
(	2205	)	,
(	2201	)	,
(	2196	)	,
(	2192	)	,
(	2188	)	,
(	2184	)	,
(	2180	)	,
(	2176	)	,
(	2172	)	,
(	2168	)	,
(	2164	)	,
(	2160	)	,
(	2156	)	,
(	2152	)	,
(	2148	)	,
(	2144	)	,
(	2140	)	,
(	2136	)	,
(	2132	)	,
(	2128	)	,
(	2124	)	,
(	2120	)	,
(	2117	)	,
(	2113	)	,
(	2109	)	,
(	2105	)	,
(	2101	)	,
(	2097	)	,
(	2093	)	,
(	2090	)	,
(	2086	)	,
(	2082	)	,
(	2078	)	,
(	2075	)	,
(	2071	)	,
(	2067	)	,
(	2063	)	,
(	2060	)	,
(	2056	)	,
(	2052	)	,
(	2049	)	,
(	2045	)	,
(	2041	)	,
(	2038	)	,
(	2034	)	,
(	2030	)	,
(	2027	)	,
(	2023	)	,
(	2020	)	,
(	2016	)	,
(	2012	)	,
(	2009	)	,
(	2005	)	,
(	2002	)	,
(	1998	)	,
(	1995	)	,
(	1991	)	,
(	1988	)	,
(	1984	)	,
(	1981	)	,
(	1977	)	,
(	1974	)	,
(	1970	)	,
(	1967	)	,
(	1964	)	,
(	1960	)	,
(	1957	)	,
(	1953	)	,
(	1950	)	,
(	1947	)	,
(	1943	)	,
(	1940	)	,
(	1937	)	,
(	1933	)	,
(	1930	)	,
(	1927	)	,
(	1923	)	,
(	1920	)	,
(	1917	)	,
(	1914	)	,
(	1910	)	,
(	1907	)	,
(	1904	)	,
(	1901	)	,
(	1897	)	,
(	1894	)	,
(	1891	)	,
(	1888	)	,
(	1885	)	,
(	1881	)	,
(	1878	)	,
(	1875	)	,
(	1872	)	,
(	1869	)	,
(	1866	)	,
(	1863	)	,
(	1860	)	,
(	1856	)	,
(	1853	)	,
(	1850	)	,
(	1847	)	,
(	1844	)	,
(	1841	)	,
(	1838	)	,
(	1835	)	,
(	1832	)	,
(	1829	)	,
(	1826	)	,
(	1823	)	,
(	1820	)	,
(	1817	)	,
(	1814	)	,
(	1811	)	,
(	1808	)	,
(	1805	)	,
(	1802	)	,
(	1799	)	,
(	1797	)	,
(	1794	)	,
(	1791	)	,
(	1788	)	,
(	1785	)	,
(	1782	)	,
(	1779	)	,
(	1776	)	,
(	1774	)	,
(	1771	)	,
(	1768	)	,
(	1765	)	,
(	1762	)	,
(	1760	)	,
(	1757	)	,
(	1754	)	,
(	1751	)	,
(	1748	)	,
(	1746	)	,
(	1743	)	,
(	1740	)	,
(	1738	)	,
(	1735	)	,
(	1732	)	,
(	1729	)	,
(	1727	)	,
(	1724	)	,
(	1721	)	,
(	1719	)	,
(	1716	)	,
(	1713	)	,
(	1711	)	,
(	1708	)	,
(	1706	)	,
(	1703	)	,
(	1700	)	,
(	1698	)	,
(	1695	)	,
(	1693	)	,
(	1690	)	,
(	1687	)	,
(	1685	)	,
(	1682	)	,
(	1680	)	,
(	1677	)	,
(	1675	)	,
(	1672	)	,
(	1670	)	,
(	1667	)	,
(	1665	)	,
(	1662	)	,
(	1660	)	,
(	1657	)	,
(	1655	)	,
(	1652	)	,
(	1650	)	,
(	1647	)	,
(	1645	)	,
(	1643	)	,
(	1640	)	,
(	1638	)	,
(	1635	)	,
(	1633	)	,
(	1630	)	,
(	1628	)	,
(	1626	)	,
(	1623	)	,
(	1621	)	,
(	1619	)	,
(	1616	)	,
(	1614	)	,
(	1612	)	,
(	1609	)	,
(	1607	)	,
(	1605	)	,
(	1602	)	,
(	1600	)	,
(	1598	)	,
(	1596	)	,
(	1593	)	,
(	1591	)	,
(	1589	)	,
(	1586	)	,
(	1584	)	,
(	1582	)	,
(	1580	)	,
(	1578	)	,
(	1575	)	,
(	1573	)	,
(	1571	)	,
(	1569	)	,
(	1567	)	,
(	1564	)	,
(	1562	)	,
(	1560	)	,
(	1558	)	,
(	1556	)	,
(	1554	)	,
(	1551	)	,
(	1549	)	,
(	1547	)	,
(	1545	)	,
(	1543	)	,
(	1541	)	,
(	1539	)	,
(	1537	)	,
(	1535	)	,
(	1532	)	,
(	1530	)	,
(	1528	)	,
(	1526	)	,
(	1524	)	,
(	1522	)	,
(	1520	)	,
(	1518	)	,
(	1516	)	,
(	1514	)	,
(	1512	)	,
(	1510	)	,
(	1508	)	,
(	1506	)	,
(	1504	)	,
(	1502	)	,
(	1500	)	,
(	1498	)	,
(	1496	)	,
(	1494	)	,
(	1492	)	,
(	1490	)	,
(	1488	)	,
(	1486	)	,
(	1484	)	,
(	1482	)	,
(	1481	)	,
(	1479	)	,
(	1477	)	,
(	1475	)	,
(	1473	)	,
(	1471	)	,
(	1469	)	,
(	1467	)	,
(	1465	)	,
(	1464	)	,
(	1462	)	,
(	1460	)	,
(	1458	)	,
(	1456	)	,
(	1454	)	,
(	1453	)	,
(	1451	)	,
(	1449	)	,
(	1447	)	,
(	1445	)	,
(	1443	)	,
(	1442	)	,
(	1440	)	,
(	1438	)	,
(	1436	)	,
(	1435	)	,
(	1433	)	,
(	1431	)	,
(	1429	)	,
(	1427	)	,
(	1426	)	,
(	1424	)	,
(	1422	)	,
(	1421	)	,
(	1419	)	,
(	1417	)	,
(	1415	)	,
(	1414	)	,
(	1412	)	,
(	1410	)	,
(	1409	)	,
(	1407	)	,
(	1405	)	,
(	1404	)	,
(	1402	)	,
(	1400	)	,
(	1399	)	,
(	1397	)	,
(	1395	)	,
(	1394	)	,
(	1392	)	,
(	1390	)	,
(	1389	)	,
(	1387	)	,
(	1385	)	,
(	1384	)	,
(	1382	)	,
(	1381	)	,
(	1379	)	,
(	1377	)	,
(	1376	)	,
(	1374	)	,
(	1373	)	,
(	1371	)	,
(	1369	)	,
(	1368	)	,
(	1366	)	,
(	1365	)	,
(	1363	)	,
(	1362	)	,
(	1360	)	,
(	1359	)	,
(	1357	)	,
(	1356	)	,
(	1354	)	,
(	1352	)	,
(	1351	)	,
(	1349	)	,
(	1348	)	,
(	1346	)	,
(	1345	)	,
(	1343	)	,
(	1342	)	,
(	1340	)	,
(	1339	)	,
(	1338	)	,
(	1336	)	,
(	1335	)	,
(	1333	)	,
(	1332	)	,
(	1330	)	,
(	1329	)	,
(	1327	)	,
(	1326	)	,
(	1324	)	,
(	1323	)	,
(	1322	)	,
(	1320	)	,
(	1319	)	,
(	1317	)	,
(	1316	)	,
(	1315	)	,
(	1313	)	,
(	1312	)	,
(	1310	)	,
(	1309	)	,
(	1308	)	,
(	1306	)	,
(	1305	)	,
(	1303	)	,
(	1302	)	,
(	1301	)	,
(	1299	)	,
(	1298	)	,
(	1297	)	,
(	1295	)	,
(	1294	)	,
(	1293	)	,
(	1291	)	,
(	1290	)	,
(	1289	)	,
(	1287	)	,
(	1286	)	,
(	1285	)	,
(	1283	)	,
(	1282	)	,
(	1281	)	,
(	1279	)	,
(	1278	)	,
(	1277	)	,
(	1276	)	,
(	1274	)	,
(	1273	)	,
(	1272	)	,
(	1270	)	,
(	1269	)	,
(	1268	)	,
(	1267	)	,
(	1265	)	,
(	1264	)	,
(	1263	)	,
(	1262	)	,
(	1260	)	,
(	1259	)	,
(	1258	)	,
(	1257	)	,
(	1255	)	,
(	1254	)	,
(	1253	)	,
(	1252	)	,
(	1251	)	,
(	1249	)	,
(	1248	)	,
(	1247	)	,
(	1246	)	,
(	1244	)	,
(	1243	)	,
(	1242	)	,
(	1241	)	,
(	1240	)	,
(	1239	)	,
(	1237	)	,
(	1236	)	,
(	1235	)	,
(	1234	)	,
(	1233	)	,
(	1232	)	,
(	1230	)	,
(	1229	)	,
(	1228	)	,
(	1227	)	,
(	1226	)	,
(	1225	)	,
(	1223	)	,
(	1222	)	,
(	1221	)	,
(	1220	)	,
(	1219	)	,
(	1218	)	,
(	1217	)	,
(	1216	)	,
(	1214	)	,
(	1213	)	,
(	1212	)	,
(	1211	)	,
(	1210	)	,
(	1209	)	,
(	1208	)	,
(	1207	)	,
(	1206	)	,
(	1205	)	,
(	1203	)	,
(	1202	)	,
(	1201	)	,
(	1200	)	,
(	1199	)	,
(	1198	)	,
(	1197	)	,
(	1196	)	,
(	1195	)	,
(	1194	)	,
(	1193	)	,
(	1192	)	,
(	1191	)	,
(	1190	)	,
(	1189	)	,
(	1188	)	,
(	1187	)	,
(	1186	)	,
(	1184	)	,
(	1183	)	,
(	1182	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1178	)	,
(	1177	)	,
(	1176	)	,
(	1175	)	,
(	1174	)	,
(	1173	)	,
(	1172	)	,
(	1171	)	,
(	1170	)	,
(	1169	)	,
(	1168	)	,
(	1167	)	,
(	1166	)	,
(	1165	)	,
(	1164	)	,
(	1163	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1159	)	,
(	1159	)	,
(	1158	)	,
(	1157	)	,
(	1156	)	,
(	1155	)	,
(	1154	)	,
(	1153	)	,
(	1152	)	,
(	1151	)	,
(	1150	)	,
(	1149	)	,
(	1148	)	,
(	1147	)	,
(	1146	)	,
(	1145	)	,
(	1144	)	,
(	1143	)	,
(	1142	)	,
(	1142	)	,
(	1141	)	,
(	1140	)	,
(	1139	)	,
(	1138	)	,
(	1137	)	,
(	1136	)	,
(	1135	)	,
(	1134	)	,
(	1133	)	,
(	1132	)	,
(	1132	)	,
(	1131	)	,
(	1130	)	,
(	1129	)	,
(	1128	)	,
(	1127	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1121	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1117	)	,
(	1116	)	,
(	1115	)	,
(	1114	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1105	)	,
(	1105	)	,
(	1104	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1100	)	,
(	1099	)	,
(	1098	)	,
(	1097	)	,
(	1096	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1091	)	,
(	1090	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1083	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1080	)	,
(	1079	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1069	)	,
(	1068	)	,
(	1067	)	,
(	1066	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1054	)	,
(	1053	)	,
(	1052	)	,
(	1051	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1048	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1031	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1026	)	,
(	1025	)	,
(	1024	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1019	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1007	)	,
(	1006	)	,
(	1005	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1001	)	,
(	1000	)	,
(	999	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	991	)	,
(	990	)	,
(	990	)	,
(	989	)	,
(	988	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	986	)	,
(	985	)	,
(	984	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	980	)	,
(	979	)	,
(	979	)	,
(	978	)	,
(	977	)	,
(	977	)	,
(	976	)	,
(	975	)	,
(	975	)	,
(	974	)	,
(	974	)	,
(	973	)	,
(	972	)	,
(	972	)	,
(	971	)	,
(	970	)	,
(	970	)	,
(	969	)	,
(	968	)	,
(	968	)	,
(	967	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	963	)	,
(	962	)	,
(	962	)	,
(	961	)	,
(	960	)	,
(	960	)	,
(	959	)	,
(	958	)	,
(	958	)	,
(	957	)	,
(	957	)	,
(	956	)	,
(	955	)	,
(	955	)	,
(	954	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	952	)	,
(	951	)	,
(	950	)	,
(	950	)	,
(	949	)	,
(	949	)	,
(	948	)	,
(	947	)	,
(	947	)	,
(	946	)	,
(	946	)	,
(	945	)	,
(	944	)	,
(	944	)	,
(	943	)	,
(	943	)	,
(	942	)	,
(	941	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	939	)	,
(	938	)	,
(	938	)	,
(	937	)	,
(	936	)	,
(	936	)	,
(	935	)	,
(	935	)	,
(	934	)	,
(	933	)	,
(	933	)	,
(	932	)	,
(	932	)	,
(	931	)	,
(	930	)	,
(	930	)	,
(	929	)	,
(	929	)	,
(	928	)	,
(	927	)	,
(	927	)	,
(	926	)	,
(	926	)	,
(	925	)	,
(	924	)	,
(	924	)	,
(	923	)	,
(	923	)	,
(	922	)	,
(	921	)	,
(	921	)	,
(	920	)	,
(	920	)	,
(	919	)	,
(	918	)	,
(	918	)	,
(	917	)	,
(	917	)	,
(	916	)	,
(	915	)	,
(	915	)	,
(	914	)	,
(	914	)	,
(	913	)	,
(	912	)	,
(	912	)	,
(	911	)	,
(	911	)	,
(	910	)	,
(	909	)	,
(	909	)	,
(	908	)	,
(	908	)	,
(	907	)	,
(	907	)	,
(	906	)	,
(	905	)	,
(	905	)	,
(	904	)	,
(	904	)	,
(	903	)	,
(	902	)	,
(	902	)	,
(	901	)	,
(	901	)	,
(	900	)	,
(	899	)	,
(	899	)	,
(	898	)	,
(	898	)	,
(	897	)	,
(	896	)	,
(	896	)	,
(	895	)	,
(	895	)	,
(	894	)	,
(	894	)	,
(	893	)	,
(	892	)	,
(	892	)	,
(	891	)	,
(	891	)	,
(	890	)	,
(	889	)	,
(	889	)	,
(	888	)	,
(	888	)	,
(	887	)	,
(	886	)	,
(	886	)	,
(	885	)	,
(	885	)	,
(	884	)	,
(	884	)	,
(	883	)	,
(	882	)	,
(	882	)	,
(	881	)	,
(	881	)	,
(	880	)	,
(	879	)	,
(	879	)	,
(	878	)	,
(	878	)	,
(	877	)	,
(	877	)	,
(	876	)	,
(	875	)	,
(	875	)	,
(	874	)	,
(	874	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	868	)	,
(	868	)	,
(	867	)	,
(	867	)	,
(	866	)	,
(	865	)	,
(	865	)	,
(	864	)	,
(	864	)	,
(	863	)	,
(	863	)	,
(	862	)	,
(	861	)	,
(	861	)	,
(	860	)	,
(	860	)	,
(	859	)	,
(	858	)	,
(	858	)	,
(	857	)	,
(	857	)	,
(	856	)	,
(	856	)	,
(	855	)	,
(	854	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	851	)	,
(	851	)	,
(	850	)	,
(	850	)	,
(	849	)	,
(	849	)	,
(	848	)	,
(	847	)	,
(	847	)	,
(	846	)	,
(	846	)	,
(	845	)	,
(	845	)	,
(	844	)	,
(	843	)	,
(	843	)	,
(	842	)	,
(	842	)	,
(	841	)	,
(	840	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	838	)	,
(	837	)	,
(	836	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	834	)	,
(	833	)	,
(	832	)	,
(	832	)	,
(	831	)	,
(	831	)	,
(	830	)	,
(	829	)	,
(	829	)	,
(	828	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	824	)	,
(	823	)	,
(	823	)	,
(	822	)	,
(	821	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	817	)	,
(	816	)	,
(	816	)	,
(	815	)	,
(	814	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	812	)	,
(	811	)	,
(	810	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	807	)	,
(	807	)	,
(	806	)	,
(	806	)	,
(	805	)	,
(	805	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	797	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	794	)	,
(	793	)	,
(	792	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	782	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	769	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	761	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	759	)	,
(	758	)	,
(	757	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	755	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	748	)	,
(	747	)	,
(	747	)	,
(	746	)	,
(	746	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	742	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	738	)	,
(	737	)	,
(	736	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	730	)	,
(	729	)	,
(	728	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	719	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	716	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	699	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	697	)	,
(	696	)	,
(	696	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	683	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	679	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	672	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	667	)	,
(	666	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	664	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	655	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	647	)	,
(	646	)	,
(	646	)	,
(	645	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	643	)	,
(	642	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	639	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	617	)	,
(	616	)	,
(	616	)	,
(	615	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	608	)	,
(	607	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	596	)	,
(	595	)	,
(	595	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	592	)	,
(	591	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	574	)	,
(	573	)	,
(	573	)	,
(	572	)	,
(	572	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	567	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	564	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	559	)	,
(	558	)	,
(	558	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	551	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	548	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	540	)	,
(	539	)	,
(	539	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	537	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	399	)	,
(	398	)	,
(	398	)	,
(	397	)	,
(	397	)	,
(	396	)	,
(	396	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	393	)	,
(	393	)	,
(	392	)	,
(	392	)	,
(	391	)	,
(	390	)	,
(	390	)	,
(	389	)	,
(	389	)	,
(	388	)	,
(	387	)	,
(	387	)	,
(	386	)	,
(	386	)	,
(	385	)	,
(	384	)	,
(	384	)	,
(	383	)	,
(	382	)	,
(	382	)	,
(	381	)	,
(	380	)	,
(	380	)	,
(	379	)	,
(	378	)	,
(	378	)	,
(	377	)	,
(	376	)	,
(	376	)	,
(	375	)	,
(	374	)	,
(	374	)	,
(	373	)	,
(	372	)	,
(	372	)	,
(	371	)	,
(	370	)	,
(	369	)	,
(	369	)	,
(	368	)	,
(	367	)	,
(	367	)	,
(	366	)	,
(	365	)	,
(	364	)	,
(	364	)	,
(	363	)	,
(	362	)	,
(	361	)	,
(	360	)	,
(	360	)	,
(	359	)	,
(	358	)	,
(	357	)	,
(	357	)	,
(	356	)	,
(	355	)	,
(	354	)	,
(	353	)	,
(	353	)	,
(	352	)	,
(	351	)	,
(	350	)	,
(	349	)	,
(	348	)	,
(	347	)	,
(	347	)	,
(	346	)	,
(	345	)	,
(	344	)	,
(	343	)	,
(	342	)	,
(	341	)	,
(	341	)	,
(	340	)	,
(	339	)	,
(	338	)	,
(	337	)	,
(	336	)	,
(	335	)	,
(	334	)	,
(	333	)	,
(	332	)	,
(	331	)	,
(	330	)	,
(	329	)	,
(	329	)	,
(	328	)	,
(	327	)	,
(	326	)	,
(	325	)	,
(	324	)	,
(	323	)	,
(	322	)	,
(	321	)	,
(	320	)	,
(	319	)	,
(	318	)	,
(	317	)	,
(	316	)	,
(	315	)	,
(	314	)	,
(	313	)	,
(	311	)	,
(	310	)	,
(	309	)	,
(	308	)	,
(	307	)	,
(	306	)	,
(	305	)	,
(	304	)	,
(	303	)	,
(	302	)	,
(	301	)	,
(	300	)	,
(	298	)	,
(	297	)	,
(	296	)	,
(	295	)	,
(	294	)	,
(	293	)	,
(	292	)	,
(	290	)	,
(	289	)	,
(	288	)	,
(	287	)	,
(	286	)	,
(	285	)	,
(	283	)	,
(	282	)	,
(	281	)	,
(	280	)	,
(	279	)	,
(	277	)	,
(	276	)	,
(	275	)	,
(	274	)	,
(	272	)	,
(	271	)	,
(	270	)	,
(	269	)	,
(	267	)	,
(	266	)	,
(	265	)	,
(	263	)	,
(	262	)	,
(	261	)	,
(	259	)	,
(	258	)	,
(	257	)	,
(	255	)	,
(	254	)	,
(	253	)	,
(	251	)	,
(	250	)	,
(	249	)	,
(	247	)	,
(	246	)	,
(	245	)	,
(	243	)	,
(	242	)	,
(	240	)	,
(	239	)	,
(	237	)	,
(	236	)	,
(	235	)	,
(	233	)	,
(	232	)	,
(	230	)	,
(	229	)	,
(	227	)	,
(	226	)	,
(	224	)	,
(	223	)	,
(	221	)	,
(	220	)	,
(	218	)	,
(	217	)	,
(	215	)	,
(	214	)	,
(	212	)	,
(	211	)	,
(	209	)	,
(	207	)	,
(	206	)	,
(	204	)	,
(	203	)	,
(	201	)	,
(	200	)	,
(	198	)	,
(	196	)	,
(	195	)	,
(	193	)	,
(	191	)	,
(	190	)	,
(	188	)	,
(	186	)	,
(	185	)	,
(	183	)	,
(	181	)	,
(	180	)	,
(	178	)	,
(	176	)	,
(	175	)	,
(	173	)	,
(	171	)	,
(	169	)	,
(	168	)	,
(	166	)	,
(	164	)	,
(	162	)	,
(	160	)	,
(	159	)	,
(	157	)	,
(	155	)	,
(	153	)	,
(	151	)	,
(	150	)	,
(	148	)	,
(	146	)	,
(	144	)	,
(	142	)	,
(	140	)	,
(	138	)	,
(	136	)	,
(	135	)	,
(	133	)	,
(	131	)	,
(	129	)	,
(	127	)	,
(	125	)	,
(	123	)	,
(	121	)	,
(	119	)	,
(	117	)	,
(	115	)	,
(	113	)	,
(	111	)	,
(	109	)	,
(	107	)	,
(	105	)	,
(	103	)	,
(	101	)	,
(	99	)	,
(	97	)	,
(	95	)	,
(	93	)	,
(	90	)	,
(	88	)	,
(	86	)	,
(	84	)	,
(	82	)	,
(	80	)	,
(	78	)	,
(	76	)	,
(	73	)	,
(	71	)	,
(	69	)	,
(	67	)	,
(	65	)	,
(	62	)	,
(	60	)	,
(	58	)	,
(	56	)	,
(	53	)	,
(	51	)	,
(	49	)	,
(	47	)	,
(	44	)	,
(	42	)	,
(	40	)	,
(	37	)	,
(	35	)	,
(	33	)	,
(	30	)	,
(	28	)	,
(	26	)	,
(	23	)	,
(	21	)	,
(	18	)	,
(	16	)	,
(	14	)	,
(	11	)	,
(	9	)	,
(	6	)	,
(	4	)	,
(	1	)	,
(	-1	)	,
(	-4	)	,
(	-6	)	,
(	-9	)	,
(	-11	)	,
(	-14	)	,
(	-16	)	,
(	-19	)	,
(	-21	)	,
(	-24	)	,
(	-27	)	,
(	-29	)	,
(	-32	)	,
(	-34	)	,
(	-37	)	,
(	-40	)	,
(	-42	)	,
(	-45	)	,
(	-48	)	,
(	-50	)	,
(	-53	)	,
(	-56	)	,
(	-58	)	,
(	-61	)	,
(	-64	)	,
(	-67	)	,
(	-69	)	,
(	-72	)	,
(	-75	)	,
(	-78	)	,
(	-81	)	,
(	-83	)	,
(	-86	)	,
(	-89	)	,
(	-92	)	,
(	-95	)	,
(	-98	)	,
(	-100	)	,
(	-103	)	,
(	-106	)	,
(	-109	)	,
(	-112	)	,
(	-115	)	,
(	-118	)	,
(	-121	)	,
(	-124	)	,
(	-127	)	,
(	-130	)	,
(	-133	)	,
(	-136	)	,
(	-139	)	,
(	-142	)	,
(	-145	)	,
(	-148	)	,
(	-151	)	,
(	-154	)	,
(	-157	)	,
(	-161	)	,
(	-164	)	,
(	-167	)	,
(	-170	)	,
(	-173	)	,
(	-176	)	,
(	-179	)	,
(	-183	)	,
(	-186	)	,
(	-189	)	,
(	-192	)	,
(	-196	)	,
(	-199	)	,
(	-202	)	,
(	-205	)	,
(	-209	)	,
(	-212	)	,
(	-215	)	,
(	-219	)	,
(	-222	)	,
(	-225	)	,
(	-229	)	,
(	-232	)	,
(	-236	)	,
(	-239	)	,
(	-242	)	,
(	-246	)	,
(	-249	)	,
(	-253	)	,
(	-256	)	,
(	-260	)	,
(	-263	)	,
(	-267	)	,
(	-270	)	,
(	-274	)	,
(	-277	)	,
(	-281	)	,
(	-284	)	,
(	-288	)	,
(	-292	)	,
(	-295	)	,
(	-299	)	,
(	-303	)	,
(	-306	)	,
(	-310	)	,
(	-314	)	,
(	-317	)	,
(	-321	)	,
(	-325	)	,
(	-328	)	,
(	-332	)	,
(	-336	)	,
(	-340	)	,
(	-344	)	,
(	-347	)	,
(	-351	)	,
(	-355	)	,
(	-359	)	,
(	-363	)	,
(	-367	)	,
(	-370	)	,
(	-374	)	,
(	-378	)	,
(	-382	)	,
(	-386	)	,
(	-390	)	,
(	-394	)	,
(	-398	)	,
(	-402	)	,
(	-406	)	,
(	-410	)	,
(	-414	)	,
(	-418	)	,
(	-422	)	,
(	-426	)	,
(	-431	)	,
(	-435	)	,
(	-439	)	,
(	-443	)	,
(	-447	)	,
(	-451	)	,
(	-455	)	,
(	-460	)	,
(	-464	)	,
(	-468	)	,
(	-472	)	,
(	-477	)	,
(	-481	)	,
(	-485	)	,
(	-490	)	,
(	-494	)	,
(	-498	)	,
(	-503	)	,
(	-507	)	,
(	-511	)	,
(	-516	)	,
(	-520	)	,
(	-525	)	,
(	-529	)	,
(	-533	)	,
(	-538	)	,
(	-542	)	,
(	-547	)	,
(	-551	)	,
(	-556	)	,
(	-561	)	,
(	-565	)	,
(	-570	)	,
(	-574	)	,
(	-579	)	,
(	-584	)	,
(	-588	)	,
(	-593	)	,
(	-598	)	,
(	-602	)	,
(	-607	)	,
(	-612	)	,
(	-617	)	,
(	-621	)	,
(	-626	)	,
(	-631	)	,
(	-636	)	,
(	-640	)	,
(	-645	)	,
(	-650	)	,
(	-655	)	,
(	-660	)	,
(	-665	)	,
(	-670	)	,
(	-675	)	,
(	-680	)	,
(	-685	)	,
(	-690	)	,
(	-695	)	,
(	-700	)	,
(	-705	)	,
(	-710	)	,
(	-715	)	,
(	-720	)	,
(	-725	)	,
(	-730	)	,
(	-735	)	,
(	-741	)	,
(	-746	)	,
(	-751	)	,
(	-756	)	,
(	-761	)	,
(	-767	)	,
(	-772	)	,
(	-777	)	,
(	-782	)	,
(	-788	)	,
(	-793	)	,
(	-798	)	,
(	-804	)	,
(	-809	)	,
(	-815	)	,
(	-820	)	,
(	-825	)	,
(	-831	)	,
(	-836	)	,
(	-842	)	,
(	-847	)	,
(	-853	)	,
(	-858	)	,
(	-864	)	,
(	-870	)	,
(	-875	)	,
(	-881	)	,
(	-886	)	,
(	-892	)	,
(	-898	)	,
(	-903	)	,
(	-909	)	,
(	-915	)	,
(	-921	)	,
(	-926	)	,
(	-932	)	,
(	-938	)	,
(	-944	)	,
(	-950	)	,
(	-955	)	,
(	-961	)	,
(	-967	)	,
(	-973	)	,
(	-979	)	,
(	-985	)	,
(	-991	)	,
(	-997	)	,
(	-1003	)	,
(	-1009	)	,
(	-1015	)	,
(	-1021	)	,
(	-1027	)	,
(	-1033	)	,
(	-1039	)	,
(	-1046	)	,
(	-1052	)	,
(	-1058	)	,
(	-1064	)	,
(	-1070	)	,
(	-1077	)	,
(	-1083	)	,
(	-1089	)	,
(	-1095	)	,
(	-1102	)	,
(	-1108	)	,
(	-1114	)	,
(	-1121	)	,
(	-1127	)	,
(	-1134	)	,
(	-1140	)	,
(	-1146	)	,
(	-1153	)	,
(	-1159	)	,
(	-1166	)	,
(	-1172	)	,
(	-1179	)	,
(	-1186	)	,
(	-1192	)	,
(	-1199	)	,
(	-1205	)	,
(	-1212	)	,
(	-1219	)	,
(	-1225	)	,
(	-1232	)	,
(	-1239	)	,
(	-1246	)	,
(	-1252	)	,
(	-1259	)	,
(	-1266	)	,
(	-1273	)	,
(	-1280	)	,
(	-1287	)	,
(	-1294	)	,
(	-1301	)	,
(	-1307	)	,
(	-1314	)	,
(	-1321	)	,
(	-1328	)	,
(	-1335	)	,
(	-1343	)	,
(	-1350	)	,
(	-1357	)	,
(	-1364	)	,
(	-1371	)	,
(	-1378	)	,
(	-1385	)	,
(	-1392	)	,
(	-1400	)	,
(	-1407	)	,
(	-1414	)	,
(	-1421	)	,
(	-1429	)	,
(	-1436	)	,
(	-1443	)	,
(	-1451	)	,
(	-1458	)	,
(	-1466	)	,
(	-1473	)	,
(	-1481	)	,
(	-1488	)	,
(	-1496	)	,
(	-1503	)	,
(	-1511	)	,
(	-1518	)	,
(	-1526	)	,
(	-1533	)	,
(	-1541	)	,
(	-1549	)	,
(	-1556	)	,
(	-1564	)	,
(	-1572	)	,
(	-1580	)	,
(	-1587	)	,
(	-1595	)	,
(	-1603	)	,
(	-1611	)	,
(	-1619	)	,
(	-1627	)	,
(	-1635	)	,
(	-1642	)	,
(	-1650	)	,
(	-1658	)	,
(	-1666	)	,
(	-1674	)	,
(	-1683	)	,
(	-1691	)	,
(	-1699	)	,
(	-1707	)	,
(	-1715	)	,
(	-1723	)	,
(	-1731	)	,
(	-1740	)	,
(	-1748	)	,
(	-1756	)	,
(	-1764	)	,
(	-1773	)	,
(	-1781	)	,
(	-1789	)	,
(	-1798	)	,
(	-1806	)	,
(	-1815	)	,
(	-1823	)	,
(	-1832	)	,
(	-1840	)	,
(	-1849	)	,
(	-1857	)	,
(	-1866	)	,
(	-1874	)	,
(	-1883	)	,
(	-1892	)	,
(	-1900	)	,
(	-1909	)	,
(	-1918	)	,
(	-1926	)	,
(	-1935	)	,
(	-1944	)	,
(	-1953	)	,
(	-1962	)	,
(	-1971	)	,
(	-1980	)	,
(	-1988	)	,
(	-1997	)	,
(	-2006	)	,
(	-2015	)	,
(	-2024	)	,
(	-2033	)	,
(	-2043	)	,
(	-2052	)	,
(	-2061	)	,
(	-2070	)	,
(	-2079	)	,
(	-2088	)	,
(	-2098	)	,
(	-2107	)	,
(	-2116	)	,
(	-2125	)	,
(	-2135	)	,
(	-2144	)	,
(	-2153	)	,
(	-2163	)	,
(	-2172	)	,
(	-2182	)	,
(	-2191	)	,
(	-2201	)	,
(	-2210	)	,
(	-2220	)	,
(	-2230	)	,
(	-2239	)	,
(	-2249	)	,
(	-2258	)	,
(	-2268	)	,
(	-2278	)	,
(	-2288	)	,
(	-2297	)	,
(	-2307	)	,
(	-2317	)	,
(	-2327	)	,
(	-2337	)	,
(	-2347	)	,
(	-2357	)	,
(	-2367	)	,
(	-2377	)	,
(	-2387	)	,
(	-2397	)	,
(	-2407	)	,
(	-2417	)	,
(	-2427	)	,
(	-2437	)	,
(	-2447	)	,
(	-2458	)	,
(	-2468	)	,
(	-2478	)	,
(	-2489	)	,
(	-2499	)	,
(	-2509	)	,
(	-2520	)	,
(	-2530	)	,
(	-2540	)	,
(	-2551	)	,
(	-2561	)	,
(	-2572	)	,
(	-2583	)	,
(	-2593	)	,
(	-2604	)	,
(	-2614	)	,
(	-2625	)	,
(	-2636	)	,
(	-2646	)	,
(	-2657	)	,
(	-2668	)	,
(	-2679	)	,
(	-2690	)	,
(	-2701	)	,
(	-2711	)	,
(	-2722	)	,
(	-2733	)	,
(	-2744	)	,
(	-2755	)	,
(	-2766	)	,
(	-2777	)	,
(	-2789	)	,
(	-2800	)	,
(	-2811	)	,
(	-2822	)	,
(	-2833	)	,
(	-2844	)	,
(	-2856	)	,
(	-2867	)	,
(	-2878	)	,
(	-2890	)	,
(	-2901	)	,
(	-2913	)	,
(	-2924	)	,
(	-2936	)	,
(	-2947	)	,
(	-2959	)	,
(	-2970	)	,
(	-2982	)	,
(	-2993	)	,
(	-3005	)	,
(	-3017	)	,
(	-3029	)	,
(	-3040	)	,
(	-3052	)	,
(	-3064	)	,
(	-3076	)	,
(	-3088	)	,
(	-3100	)	,
(	-3112	)	,
(	-3124	)	,
(	-3136	)	,
(	-3148	)	,
(	-3160	)	,
(	-3172	)	,
(	-3184	)	,
(	-3196	)	,
(	-3208	)	,
(	-3221	)	,
(	-3233	)	,
(	-3245	)	,
(	-3257	)	,
(	-3270	)	,
(	-3282	)	,
(	-3295	)	,
(	-3307	)	,
(	-3320	)	,
(	-3332	)	,
(	-3345	)	,
(	-3357	)	,
(	-3370	)	,
(	-3382	)	,
(	-3395	)	,
(	-3408	)	,
(	-3421	)	,
(	-3433	)	,
(	-3446	)	,
(	-3459	)	,
(	-3472	)	,
(	-3485	)	,
(	-3498	)	,
(	-3511	)	,
(	-3524	)	,
(	-3537	)	,
(	-3550	)	,
(	-3563	)	,
(	-3576	)	,
(	-3589	)	,
(	-3602	)	,
(	-3616	)	,
(	-3629	)	,
(	-3642	)	,
(	-3655	)	,
(	-3669	)	,
(	-3682	)	,
(	-3696	)	,
(	-3709	)	,
(	-3723	)	,
(	-3736	)	,
(	-3750	)	,
(	-3763	)	,
(	-3777	)	,
(	-3791	)	,
(	-3804	)	,
(	-3818	)	,
(	-3832	)	,
(	-3846	)	,
(	-3860	)	,
(	-3873	)	,
(	-3887	)	,
(	-3901	)	,
(	-3915	)	,
(	-3929	)	,
(	-3943	)	,
(	-3957	)	,
(	-3972	)	,
(	-3986	)	,
(	-4000	)	,
(	-4014	)	,
(	-4028	)	,
(	-4043	)	,
(	-4057	)	,
(	-4071	)	,
(	-4086	)	,
(	-4100	)	,
(	-4115	)	,
(	-4129	)	,
(	-4144	)	,
(	-4158	)	,
(	-4173	)	,
(	-4188	)	,
(	-4202	)	,
(	-4217	)	,
(	-4232	)	,
(	-4247	)	,
(	-4261	)	,
(	-4276	)	,
(	-4291	)	,
(	-4306	)	,
(	-4321	)	,
(	-4336	)	,
(	-4351	)	,
(	-4366	)	,
(	-4381	)	,
(	-4396	)	,
(	-4412	)	,
(	-4427	)	,
(	-4442	)	,
(	-4457	)	,
(	-4473	)	,
(	-4488	)	,
(	-4504	)	,
(	-4519	)	,
(	-4535	)	,
(	-4550	)	,
(	-4566	)	,
(	-4581	)	,
(	-4597	)	,
(	-4613	)	,
(	-4628	)	,
(	-4644	)	,
(	-4660	)	,
(	-4676	)	,
(	-4692	)	,
(	-4707	)	,
(	-4723	)	,
(	-4739	)	,
(	-4755	)	,
(	-4771	)	,
(	-4788	)	,
(	-4804	)	,
(	-4820	)	,
(	-4836	)	,
(	-4852	)	,
(	-4869	)	,
(	-4885	)	,
(	-4901	)	,
(	-4918	)	,
(	-4934	)	,
(	-4951	)	,
(	-4967	)	,
(	-4984	)	,
(	-5000	)	,
(	-5017	)	,
(	-5034	)	,
(	-5050	)	,
(	-5067	)	,
(	-5084	)	,
(	-5101	)	,
(	-5118	)	,
(	-5135	)	,
(	-5151	)	,
(	-5168	)	,
(	-5186	)	,
(	-5203	)	,
(	-5220	)	,
(	-5237	)	,
(	-5254	)	,
(	-5271	)	,
(	-5289	)	,
(	-5306	)	,
(	-5323	)	,
(	-5341	)	,
(	-5358	)	,
(	-5376	)	,
(	-5393	)	,
(	-5411	)	,
(	-5428	)	,
(	-5446	)	,
(	-5464	)	,
(	-5481	)	,
(	-5499	)	,
(	-5517	)	,
(	-5535	)	,
(	-5553	)	,
(	-5571	)	,
(	-5589	)	,
(	-5607	)	,
(	-5625	)	,
(	-5643	)	,
(	-5661	)	,
(	-5679	)	,
(	-5697	)	,
(	-5716	)	,
(	-5734	)	,
(	-5752	)	,
(	-5771	)	,
(	-5789	)	,
(	-5807	)	,
(	-5826	)	,
(	-5845	)	,
(	-5863	)	,
(	-5882	)	,
(	-5900	)	,
(	-5919	)	,
(	-5938	)	,
(	-5957	)	,
(	-5976	)	,
(	-5995	)	,
(	-6014	)	,
(	-6033	)	,
(	-6052	)	,
(	-6071	)	,
(	-6090	)	,
(	-6109	)	,
(	-6128	)	,
(	-6147	)	,
(	-6167	)	,
(	-6186	)	,
(	-6205	)	,
(	-6225	)	,
(	-6244	)	,
(	-6264	)	,
(	-6283	)	,
(	-6303	)	,
(	-6323	)	,
(	-6342	)	,
(	-6362	)	,
(	-6382	)	,
(	-6402	)	,
(	-6422	)	,
(	-6441	)	,
(	-6461	)	,
(	-6481	)	,
(	-6501	)	,
(	-6522	)	,
(	-6542	)	,
(	-6562	)	,
(	-6582	)	,
(	-6602	)	,
(	-6623	)	,
(	-6643	)	,
(	-6663	)	,
(	-6684	)	,
(	-6704	)	,
(	-6725	)	,
(	-6746	)	,
(	-6766	)	,
(	-6787	)	,
(	-6808	)	,
(	-6828	)	,
(	-6849	)	,
(	-6870	)	,
(	-6891	)	,
(	-6912	)	,
(	-6933	)	,
(	-6954	)	,
(	-6975	)	,
(	-6996	)	,
(	-7017	)	,
(	-7039	)	,
(	-7060	)	,
(	-7081	)	,
(	-7103	)	,
(	-7124	)	,
(	-7146	)	,
(	-7167	)	,
(	-7189	)	,
(	-7210	)	,
(	-7232	)	,
(	-7254	)	,
(	-7275	)	,
(	-7297	)	,
(	-7319	)	,
(	-7341	)	,
(	-7363	)	,
(	-7385	)	,
(	-7407	)	,
(	-7429	)	,
(	-7451	)	,
(	-7473	)	,
(	-7496	)	,
(	-7518	)	,
(	-7540	)	,
(	-7563	)	,
(	-7585	)	,
(	-7608	)	,
(	-7630	)	,
(	-7653	)	,
(	-7675	)	,
(	-7698	)	,
(	-7721	)	,
(	-7744	)	,
(	-7766	)	,
(	-7789	)	,
(	-7812	)	,
(	-7835	)	,
(	-7858	)	,
(	-7881	)	,
(	-7904	)	,
(	-7928	)	,
(	-7951	)	,
(	-7974	)	,
(	-7997	)	,
(	-8021	)	,
(	-8044	)	,
(	-8068	)	,
(	-8091	)	,
(	-8115	)	,
(	-8138	)	,
(	-8162	)	,
(	-8186	)	,
(	-8210	)	,
(	-8233	)	,
(	-8257	)	,
(	-8281	)	,
(	-8305	)	,
(	-8329	)	,
(	-8353	)	,
(	-8377	)	,
(	-8402	)	,
(	-8426	)	,
(	-8450	)	,
(	-8475	)	,
(	-8499	)	,
(	-8523	)	,
(	-8548	)	,
(	-8572	)	,
(	-8597	)	,
(	-8622	)	,
(	-8646	)	,
(	-8671	)	,
(	-8696	)	,
(	-8721	)	,
(	-8746	)	,
(	-8771	)	,
(	-8796	)	,
(	-8821	)	,
(	-8846	)	,
(	-8871	)	,
(	-8896	)	,
(	-8922	)	,
(	-8947	)	,
(	-8972	)	,
(	-8998	)	,
(	-9023	)	,
(	-9049	)	,
(	-9075	)	,
(	-9100	)	,
(	-9126	)	,
(	-9152	)	,
(	-9178	)	,
(	-9203	)	,
(	-9229	)	,
(	-9255	)	,
(	-9281	)	,
(	-9307	)	,
(	-9334	)	,
(	-9360	)	,
(	-9386	)	,
(	-9412	)	,
(	-9439	)	,
(	-9465	)	,
(	-9492	)	,
(	-9518	)	,
(	-9545	)	,
(	-9571	)	,
(	-9598	)	,
(	-9625	)	,
(	-9652	)	,
(	-9679	)	,
(	-9705	)	,
(	-9732	)	,
(	-9759	)	,
(	-9787	)	,
(	-9814	)	,
(	-9841	)	,
(	-9868	)	,
(	-9895	)	,
(	-9923	)	,
(	-9950	)	,
(	-9978	)	,
(	-10005	)	,
(	-10033	)	,
(	-10061	)	,
(	-10088	)	,
(	-10116	)	,
(	-10144	)	,
(	-10172	)	,
(	-10200	)	,
(	-10228	)	,
(	-10256	)	,
(	-10284	)	,
(	-10312	)	,
(	-10340	)	,
(	-10368	)	,
(	-10397	)	,
(	-10425	)	,
(	-10454	)	,
(	-10482	)	,
(	-10511	)	,
(	-10539	)	,
(	-10568	)	,
(	-10597	)	,
(	-10626	)	,
(	-10654	)	,
(	-10683	)	,
(	-10712	)	,
(	-10741	)	,
(	-10771	)	,
(	-10800	)	,
(	-10829	)	,
(	-10858	)	,
(	-10887	)	,
(	-10917	)	,
(	-10946	)	,
(	-10976	)	,
(	-11005	)	,
(	-11035	)	,
(	-11065	)	,
(	-11094	)	,
(	-11124	)	,
(	-11154	)	,
(	-11184	)	,
(	-11214	)	,
(	-11244	)	,
(	-11274	)	,
(	-11304	)	,
(	-11335	)	,
(	-11365	)	,
(	-11395	)	,
(	-11426	)	,
(	-11456	)	-- array index 4095 (voltage = "111111111111" or 4095 mV), distance output 3787 (37.87 cm)
);


begin
   -- This is the only statement required. It looks up the converted value of 
	-- the voltage input (in mV) in the v2d_LUT look-up table, and outputs the 
	-- distance (in 10^-4 m) in std_logic_vector format.
	process(voltage, mux_bit_close)
		begin
		if (mux_bit_close = '1') then
			distance <= std_logic_vector(to_unsigned(v2d_close(to_integer(unsigned(voltage))),distance'length));
		else
			distance <= std_logic_vector(to_unsigned(v2d_LUT(to_integer(unsigned(voltage))),distance'length));	
		end if;
	end process;

end behavior;
