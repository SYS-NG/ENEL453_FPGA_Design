LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY buzzer IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;		                         
      distance       :  IN    STD_LOGIC_VECTOR(12 DOWNTO 0);
		dac_out        :  OUT   STD_LOGIC
		);
END buzzer;

ARCHITECTURE behavior OF buzzer IS

signal counter       : unsigned(17 DOWNTO 0) := (others=>'0');
signal counter_limit : unsigned(17 DOWNTO 0);

type array_1d is array (0 to 3300) of integer;
	
constant d2count: array_1d := (
(	20000	 ),
(	20024	 ),
(	20048	 ),
(	20073	 ),
(	20097	 ),
(	20121	 ),
(	20145	 ),
(	20170	 ),
(	20194	 ),
(	20218	 ),
(	20242	 ),
(	20267	 ),
(	20291	 ),
(	20315	 ),
(	20339	 ),
(	20364	 ),
(	20388	 ),
(	20412	 ),
(	20436	 ),
(	20461	 ),
(	20485	 ),
(	20509	 ),
(	20533	 ),
(	20558	 ),
(	20582	 ),
(	20606	 ),
(	20630	 ),
(	20655	 ),
(	20679	 ),
(	20703	 ),
(	20727	 ),
(	20752	 ),
(	20776	 ),
(	20800	 ),
(	20824	 ),
(	20848	 ),
(	20873	 ),
(	20897	 ),
(	20921	 ),
(	20945	 ),
(	20970	 ),
(	20994	 ),
(	21018	 ),
(	21042	 ),
(	21067	 ),
(	21091	 ),
(	21115	 ),
(	21139	 ),
(	21164	 ),
(	21188	 ),
(	21212	 ),
(	21236	 ),
(	21261	 ),
(	21285	 ),
(	21309	 ),
(	21333	 ),
(	21358	 ),
(	21382	 ),
(	21406	 ),
(	21430	 ),
(	21455	 ),
(	21479	 ),
(	21503	 ),
(	21527	 ),
(	21552	 ),
(	21576	 ),
(	21600	 ),
(	21624	 ),
(	21648	 ),
(	21673	 ),
(	21697	 ),
(	21721	 ),
(	21745	 ),
(	21770	 ),
(	21794	 ),
(	21818	 ),
(	21842	 ),
(	21867	 ),
(	21891	 ),
(	21915	 ),
(	21939	 ),
(	21964	 ),
(	21988	 ),
(	22012	 ),
(	22036	 ),
(	22061	 ),
(	22085	 ),
(	22109	 ),
(	22133	 ),
(	22158	 ),
(	22182	 ),
(	22206	 ),
(	22230	 ),
(	22255	 ),
(	22279	 ),
(	22303	 ),
(	22327	 ),
(	22352	 ),
(	22376	 ),
(	22400	 ),
(	22424	 ),
(	22448	 ),
(	22473	 ),
(	22497	 ),
(	22521	 ),
(	22545	 ),
(	22570	 ),
(	22594	 ),
(	22618	 ),
(	22642	 ),
(	22667	 ),
(	22691	 ),
(	22715	 ),
(	22739	 ),
(	22764	 ),
(	22788	 ),
(	22812	 ),
(	22836	 ),
(	22861	 ),
(	22885	 ),
(	22909	 ),
(	22933	 ),
(	22958	 ),
(	22982	 ),
(	23006	 ),
(	23030	 ),
(	23055	 ),
(	23079	 ),
(	23103	 ),
(	23127	 ),
(	23152	 ),
(	23176	 ),
(	23200	 ),
(	23224	 ),
(	23248	 ),
(	23273	 ),
(	23297	 ),
(	23321	 ),
(	23345	 ),
(	23370	 ),
(	23394	 ),
(	23418	 ),
(	23442	 ),
(	23467	 ),
(	23491	 ),
(	23515	 ),
(	23539	 ),
(	23564	 ),
(	23588	 ),
(	23612	 ),
(	23636	 ),
(	23661	 ),
(	23685	 ),
(	23709	 ),
(	23733	 ),
(	23758	 ),
(	23782	 ),
(	23806	 ),
(	23830	 ),
(	23855	 ),
(	23879	 ),
(	23903	 ),
(	23927	 ),
(	23952	 ),
(	23976	 ),
(	24000	 ),
(	24024	 ),
(	24048	 ),
(	24073	 ),
(	24097	 ),
(	24121	 ),
(	24145	 ),
(	24170	 ),
(	24194	 ),
(	24218	 ),
(	24242	 ),
(	24267	 ),
(	24291	 ),
(	24315	 ),
(	24339	 ),
(	24364	 ),
(	24388	 ),
(	24412	 ),
(	24436	 ),
(	24461	 ),
(	24485	 ),
(	24509	 ),
(	24533	 ),
(	24558	 ),
(	24582	 ),
(	24606	 ),
(	24630	 ),
(	24655	 ),
(	24679	 ),
(	24703	 ),
(	24727	 ),
(	24752	 ),
(	24776	 ),
(	24800	 ),
(	24824	 ),
(	24848	 ),
(	24873	 ),
(	24897	 ),
(	24921	 ),
(	24945	 ),
(	24970	 ),
(	24994	 ),
(	25018	 ),
(	25042	 ),
(	25067	 ),
(	25091	 ),
(	25115	 ),
(	25139	 ),
(	25164	 ),
(	25188	 ),
(	25212	 ),
(	25236	 ),
(	25261	 ),
(	25285	 ),
(	25309	 ),
(	25333	 ),
(	25358	 ),
(	25382	 ),
(	25406	 ),
(	25430	 ),
(	25455	 ),
(	25479	 ),
(	25503	 ),
(	25527	 ),
(	25552	 ),
(	25576	 ),
(	25600	 ),
(	25624	 ),
(	25648	 ),
(	25673	 ),
(	25697	 ),
(	25721	 ),
(	25745	 ),
(	25770	 ),
(	25794	 ),
(	25818	 ),
(	25842	 ),
(	25867	 ),
(	25891	 ),
(	25915	 ),
(	25939	 ),
(	25964	 ),
(	25988	 ),
(	26012	 ),
(	26036	 ),
(	26061	 ),
(	26085	 ),
(	26109	 ),
(	26133	 ),
(	26158	 ),
(	26182	 ),
(	26206	 ),
(	26230	 ),
(	26255	 ),
(	26279	 ),
(	26303	 ),
(	26327	 ),
(	26352	 ),
(	26376	 ),
(	26400	 ),
(	26424	 ),
(	26448	 ),
(	26473	 ),
(	26497	 ),
(	26521	 ),
(	26545	 ),
(	26570	 ),
(	26594	 ),
(	26618	 ),
(	26642	 ),
(	26667	 ),
(	26691	 ),
(	26715	 ),
(	26739	 ),
(	26764	 ),
(	26788	 ),
(	26812	 ),
(	26836	 ),
(	26861	 ),
(	26885	 ),
(	26909	 ),
(	26933	 ),
(	26958	 ),
(	26982	 ),
(	27006	 ),
(	27030	 ),
(	27055	 ),
(	27079	 ),
(	27103	 ),
(	27127	 ),
(	27152	 ),
(	27176	 ),
(	27200	 ),
(	27224	 ),
(	27248	 ),
(	27273	 ),
(	27297	 ),
(	27321	 ),
(	27345	 ),
(	27370	 ),
(	27394	 ),
(	27418	 ),
(	27442	 ),
(	27467	 ),
(	27491	 ),
(	27515	 ),
(	27539	 ),
(	27564	 ),
(	27588	 ),
(	27612	 ),
(	27636	 ),
(	27661	 ),
(	27685	 ),
(	27709	 ),
(	27733	 ),
(	27758	 ),
(	27782	 ),
(	27806	 ),
(	27830	 ),
(	27855	 ),
(	27879	 ),
(	27903	 ),
(	27927	 ),
(	27952	 ),
(	27976	 ),
(	28000	 ),
(	28024	 ),
(	28048	 ),
(	28073	 ),
(	28097	 ),
(	28121	 ),
(	28145	 ),
(	28170	 ),
(	28194	 ),
(	28218	 ),
(	28242	 ),
(	28267	 ),
(	28291	 ),
(	28315	 ),
(	28339	 ),
(	28364	 ),
(	28388	 ),
(	28412	 ),
(	28436	 ),
(	28461	 ),
(	28485	 ),
(	28509	 ),
(	28533	 ),
(	28558	 ),
(	28582	 ),
(	28606	 ),
(	28630	 ),
(	28655	 ),
(	28679	 ),
(	28703	 ),
(	28727	 ),
(	28752	 ),
(	28776	 ),
(	28800	 ),
(	28824	 ),
(	28848	 ),
(	28873	 ),
(	28897	 ),
(	28921	 ),
(	28945	 ),
(	28970	 ),
(	28994	 ),
(	29018	 ),
(	29042	 ),
(	29067	 ),
(	29091	 ),
(	29115	 ),
(	29139	 ),
(	29164	 ),
(	29188	 ),
(	29212	 ),
(	29236	 ),
(	29261	 ),
(	29285	 ),
(	29309	 ),
(	29333	 ),
(	29358	 ),
(	29382	 ),
(	29406	 ),
(	29430	 ),
(	29455	 ),
(	29479	 ),
(	29503	 ),
(	29527	 ),
(	29552	 ),
(	29576	 ),
(	29600	 ),
(	29624	 ),
(	29648	 ),
(	29673	 ),
(	29697	 ),
(	29721	 ),
(	29745	 ),
(	29770	 ),
(	29794	 ),
(	29818	 ),
(	29842	 ),
(	29867	 ),
(	29891	 ),
(	29915	 ),
(	29939	 ),
(	29964	 ),
(	29988	 ),
(	30012	 ),
(	30036	 ),
(	30061	 ),
(	30085	 ),
(	30109	 ),
(	30133	 ),
(	30158	 ),
(	30182	 ),
(	30206	 ),
(	30230	 ),
(	30255	 ),
(	30279	 ),
(	30303	 ),
(	30327	 ),
(	30352	 ),
(	30376	 ),
(	30400	 ),
(	30424	 ),
(	30448	 ),
(	30473	 ),
(	30497	 ),
(	30521	 ),
(	30545	 ),
(	30570	 ),
(	30594	 ),
(	30618	 ),
(	30642	 ),
(	30667	 ),
(	30691	 ),
(	30715	 ),
(	30739	 ),
(	30764	 ),
(	30788	 ),
(	30812	 ),
(	30836	 ),
(	30861	 ),
(	30885	 ),
(	30909	 ),
(	30933	 ),
(	30958	 ),
(	30982	 ),
(	31006	 ),
(	31030	 ),
(	31055	 ),
(	31079	 ),
(	31103	 ),
(	31127	 ),
(	31152	 ),
(	31176	 ),
(	31200	 ),
(	31224	 ),
(	31248	 ),
(	31273	 ),
(	31297	 ),
(	31321	 ),
(	31345	 ),
(	31370	 ),
(	31394	 ),
(	31418	 ),
(	31442	 ),
(	31467	 ),
(	31491	 ),
(	31515	 ),
(	31539	 ),
(	31564	 ),
(	31588	 ),
(	31612	 ),
(	31636	 ),
(	31661	 ),
(	31685	 ),
(	31709	 ),
(	31733	 ),
(	31758	 ),
(	31782	 ),
(	31806	 ),
(	31830	 ),
(	31855	 ),
(	31879	 ),
(	31903	 ),
(	31927	 ),
(	31952	 ),
(	31976	 ),
(	32000	 ),
(	32024	 ),
(	32048	 ),
(	32073	 ),
(	32097	 ),
(	32121	 ),
(	32145	 ),
(	32170	 ),
(	32194	 ),
(	32218	 ),
(	32242	 ),
(	32267	 ),
(	32291	 ),
(	32315	 ),
(	32339	 ),
(	32364	 ),
(	32388	 ),
(	32412	 ),
(	32436	 ),
(	32461	 ),
(	32485	 ),
(	32509	 ),
(	32533	 ),
(	32558	 ),
(	32582	 ),
(	32606	 ),
(	32630	 ),
(	32655	 ),
(	32679	 ),
(	32703	 ),
(	32727	 ),
(	32752	 ),
(	32776	 ),
(	32800	 ),
(	32824	 ),
(	32848	 ),
(	32873	 ),
(	32897	 ),
(	32921	 ),
(	32945	 ),
(	32970	 ),
(	32994	 ),
(	33018	 ),
(	33042	 ),
(	33067	 ),
(	33091	 ),
(	33115	 ),
(	33139	 ),
(	33164	 ),
(	33188	 ),
(	33212	 ),
(	33236	 ),
(	33261	 ),
(	33285	 ),
(	33309	 ),
(	33333	 ),
(	33358	 ),
(	33382	 ),
(	33406	 ),
(	33430	 ),
(	33455	 ),
(	33479	 ),
(	33503	 ),
(	33527	 ),
(	33552	 ),
(	33576	 ),
(	33600	 ),
(	33624	 ),
(	33648	 ),
(	33673	 ),
(	33697	 ),
(	33721	 ),
(	33745	 ),
(	33770	 ),
(	33794	 ),
(	33818	 ),
(	33842	 ),
(	33867	 ),
(	33891	 ),
(	33915	 ),
(	33939	 ),
(	33964	 ),
(	33988	 ),
(	34012	 ),
(	34036	 ),
(	34061	 ),
(	34085	 ),
(	34109	 ),
(	34133	 ),
(	34158	 ),
(	34182	 ),
(	34206	 ),
(	34230	 ),
(	34255	 ),
(	34279	 ),
(	34303	 ),
(	34327	 ),
(	34352	 ),
(	34376	 ),
(	34400	 ),
(	34424	 ),
(	34448	 ),
(	34473	 ),
(	34497	 ),
(	34521	 ),
(	34545	 ),
(	34570	 ),
(	34594	 ),
(	34618	 ),
(	34642	 ),
(	34667	 ),
(	34691	 ),
(	34715	 ),
(	34739	 ),
(	34764	 ),
(	34788	 ),
(	34812	 ),
(	34836	 ),
(	34861	 ),
(	34885	 ),
(	34909	 ),
(	34933	 ),
(	34958	 ),
(	34982	 ),
(	35006	 ),
(	35030	 ),
(	35055	 ),
(	35079	 ),
(	35103	 ),
(	35127	 ),
(	35152	 ),
(	35176	 ),
(	35200	 ),
(	35224	 ),
(	35248	 ),
(	35273	 ),
(	35297	 ),
(	35321	 ),
(	35345	 ),
(	35370	 ),
(	35394	 ),
(	35418	 ),
(	35442	 ),
(	35467	 ),
(	35491	 ),
(	35515	 ),
(	35539	 ),
(	35564	 ),
(	35588	 ),
(	35612	 ),
(	35636	 ),
(	35661	 ),
(	35685	 ),
(	35709	 ),
(	35733	 ),
(	35758	 ),
(	35782	 ),
(	35806	 ),
(	35830	 ),
(	35855	 ),
(	35879	 ),
(	35903	 ),
(	35927	 ),
(	35952	 ),
(	35976	 ),
(	36000	 ),
(	36024	 ),
(	36048	 ),
(	36073	 ),
(	36097	 ),
(	36121	 ),
(	36145	 ),
(	36170	 ),
(	36194	 ),
(	36218	 ),
(	36242	 ),
(	36267	 ),
(	36291	 ),
(	36315	 ),
(	36339	 ),
(	36364	 ),
(	36388	 ),
(	36412	 ),
(	36436	 ),
(	36461	 ),
(	36485	 ),
(	36509	 ),
(	36533	 ),
(	36558	 ),
(	36582	 ),
(	36606	 ),
(	36630	 ),
(	36655	 ),
(	36679	 ),
(	36703	 ),
(	36727	 ),
(	36752	 ),
(	36776	 ),
(	36800	 ),
(	36824	 ),
(	36848	 ),
(	36873	 ),
(	36897	 ),
(	36921	 ),
(	36945	 ),
(	36970	 ),
(	36994	 ),
(	37018	 ),
(	37042	 ),
(	37067	 ),
(	37091	 ),
(	37115	 ),
(	37139	 ),
(	37164	 ),
(	37188	 ),
(	37212	 ),
(	37236	 ),
(	37261	 ),
(	37285	 ),
(	37309	 ),
(	37333	 ),
(	37358	 ),
(	37382	 ),
(	37406	 ),
(	37430	 ),
(	37455	 ),
(	37479	 ),
(	37503	 ),
(	37527	 ),
(	37552	 ),
(	37576	 ),
(	37600	 ),
(	37624	 ),
(	37648	 ),
(	37673	 ),
(	37697	 ),
(	37721	 ),
(	37745	 ),
(	37770	 ),
(	37794	 ),
(	37818	 ),
(	37842	 ),
(	37867	 ),
(	37891	 ),
(	37915	 ),
(	37939	 ),
(	37964	 ),
(	37988	 ),
(	38012	 ),
(	38036	 ),
(	38061	 ),
(	38085	 ),
(	38109	 ),
(	38133	 ),
(	38158	 ),
(	38182	 ),
(	38206	 ),
(	38230	 ),
(	38255	 ),
(	38279	 ),
(	38303	 ),
(	38327	 ),
(	38352	 ),
(	38376	 ),
(	38400	 ),
(	38424	 ),
(	38448	 ),
(	38473	 ),
(	38497	 ),
(	38521	 ),
(	38545	 ),
(	38570	 ),
(	38594	 ),
(	38618	 ),
(	38642	 ),
(	38667	 ),
(	38691	 ),
(	38715	 ),
(	38739	 ),
(	38764	 ),
(	38788	 ),
(	38812	 ),
(	38836	 ),
(	38861	 ),
(	38885	 ),
(	38909	 ),
(	38933	 ),
(	38958	 ),
(	38982	 ),
(	39006	 ),
(	39030	 ),
(	39055	 ),
(	39079	 ),
(	39103	 ),
(	39127	 ),
(	39152	 ),
(	39176	 ),
(	39200	 ),
(	39224	 ),
(	39248	 ),
(	39273	 ),
(	39297	 ),
(	39321	 ),
(	39345	 ),
(	39370	 ),
(	39394	 ),
(	39418	 ),
(	39442	 ),
(	39467	 ),
(	39491	 ),
(	39515	 ),
(	39539	 ),
(	39564	 ),
(	39588	 ),
(	39612	 ),
(	39636	 ),
(	39661	 ),
(	39685	 ),
(	39709	 ),
(	39733	 ),
(	39758	 ),
(	39782	 ),
(	39806	 ),
(	39830	 ),
(	39855	 ),
(	39879	 ),
(	39903	 ),
(	39927	 ),
(	39952	 ),
(	39976	 ),
(	40000	 ),
(	40024	 ),
(	40048	 ),
(	40073	 ),
(	40097	 ),
(	40121	 ),
(	40145	 ),
(	40170	 ),
(	40194	 ),
(	40218	 ),
(	40242	 ),
(	40267	 ),
(	40291	 ),
(	40315	 ),
(	40339	 ),
(	40364	 ),
(	40388	 ),
(	40412	 ),
(	40436	 ),
(	40461	 ),
(	40485	 ),
(	40509	 ),
(	40533	 ),
(	40558	 ),
(	40582	 ),
(	40606	 ),
(	40630	 ),
(	40655	 ),
(	40679	 ),
(	40703	 ),
(	40727	 ),
(	40752	 ),
(	40776	 ),
(	40800	 ),
(	40824	 ),
(	40848	 ),
(	40873	 ),
(	40897	 ),
(	40921	 ),
(	40945	 ),
(	40970	 ),
(	40994	 ),
(	41018	 ),
(	41042	 ),
(	41067	 ),
(	41091	 ),
(	41115	 ),
(	41139	 ),
(	41164	 ),
(	41188	 ),
(	41212	 ),
(	41236	 ),
(	41261	 ),
(	41285	 ),
(	41309	 ),
(	41333	 ),
(	41358	 ),
(	41382	 ),
(	41406	 ),
(	41430	 ),
(	41455	 ),
(	41479	 ),
(	41503	 ),
(	41527	 ),
(	41552	 ),
(	41576	 ),
(	41600	 ),
(	41624	 ),
(	41648	 ),
(	41673	 ),
(	41697	 ),
(	41721	 ),
(	41745	 ),
(	41770	 ),
(	41794	 ),
(	41818	 ),
(	41842	 ),
(	41867	 ),
(	41891	 ),
(	41915	 ),
(	41939	 ),
(	41964	 ),
(	41988	 ),
(	42012	 ),
(	42036	 ),
(	42061	 ),
(	42085	 ),
(	42109	 ),
(	42133	 ),
(	42158	 ),
(	42182	 ),
(	42206	 ),
(	42230	 ),
(	42255	 ),
(	42279	 ),
(	42303	 ),
(	42327	 ),
(	42352	 ),
(	42376	 ),
(	42400	 ),
(	42424	 ),
(	42448	 ),
(	42473	 ),
(	42497	 ),
(	42521	 ),
(	42545	 ),
(	42570	 ),
(	42594	 ),
(	42618	 ),
(	42642	 ),
(	42667	 ),
(	42691	 ),
(	42715	 ),
(	42739	 ),
(	42764	 ),
(	42788	 ),
(	42812	 ),
(	42836	 ),
(	42861	 ),
(	42885	 ),
(	42909	 ),
(	42933	 ),
(	42958	 ),
(	42982	 ),
(	43006	 ),
(	43030	 ),
(	43055	 ),
(	43079	 ),
(	43103	 ),
(	43127	 ),
(	43152	 ),
(	43176	 ),
(	43200	 ),
(	43224	 ),
(	43248	 ),
(	43273	 ),
(	43297	 ),
(	43321	 ),
(	43345	 ),
(	43370	 ),
(	43394	 ),
(	43418	 ),
(	43442	 ),
(	43467	 ),
(	43491	 ),
(	43515	 ),
(	43539	 ),
(	43564	 ),
(	43588	 ),
(	43612	 ),
(	43636	 ),
(	43661	 ),
(	43685	 ),
(	43709	 ),
(	43733	 ),
(	43758	 ),
(	43782	 ),
(	43806	 ),
(	43830	 ),
(	43855	 ),
(	43879	 ),
(	43903	 ),
(	43927	 ),
(	43952	 ),
(	43976	 ),
(	44000	 ),
(	44024	 ),
(	44048	 ),
(	44073	 ),
(	44097	 ),
(	44121	 ),
(	44145	 ),
(	44170	 ),
(	44194	 ),
(	44218	 ),
(	44242	 ),
(	44267	 ),
(	44291	 ),
(	44315	 ),
(	44339	 ),
(	44364	 ),
(	44388	 ),
(	44412	 ),
(	44436	 ),
(	44461	 ),
(	44485	 ),
(	44509	 ),
(	44533	 ),
(	44558	 ),
(	44582	 ),
(	44606	 ),
(	44630	 ),
(	44655	 ),
(	44679	 ),
(	44703	 ),
(	44727	 ),
(	44752	 ),
(	44776	 ),
(	44800	 ),
(	44824	 ),
(	44848	 ),
(	44873	 ),
(	44897	 ),
(	44921	 ),
(	44945	 ),
(	44970	 ),
(	44994	 ),
(	45018	 ),
(	45042	 ),
(	45067	 ),
(	45091	 ),
(	45115	 ),
(	45139	 ),
(	45164	 ),
(	45188	 ),
(	45212	 ),
(	45236	 ),
(	45261	 ),
(	45285	 ),
(	45309	 ),
(	45333	 ),
(	45358	 ),
(	45382	 ),
(	45406	 ),
(	45430	 ),
(	45455	 ),
(	45479	 ),
(	45503	 ),
(	45527	 ),
(	45552	 ),
(	45576	 ),
(	45600	 ),
(	45624	 ),
(	45648	 ),
(	45673	 ),
(	45697	 ),
(	45721	 ),
(	45745	 ),
(	45770	 ),
(	45794	 ),
(	45818	 ),
(	45842	 ),
(	45867	 ),
(	45891	 ),
(	45915	 ),
(	45939	 ),
(	45964	 ),
(	45988	 ),
(	46012	 ),
(	46036	 ),
(	46061	 ),
(	46085	 ),
(	46109	 ),
(	46133	 ),
(	46158	 ),
(	46182	 ),
(	46206	 ),
(	46230	 ),
(	46255	 ),
(	46279	 ),
(	46303	 ),
(	46327	 ),
(	46352	 ),
(	46376	 ),
(	46400	 ),
(	46424	 ),
(	46448	 ),
(	46473	 ),
(	46497	 ),
(	46521	 ),
(	46545	 ),
(	46570	 ),
(	46594	 ),
(	46618	 ),
(	46642	 ),
(	46667	 ),
(	46691	 ),
(	46715	 ),
(	46739	 ),
(	46764	 ),
(	46788	 ),
(	46812	 ),
(	46836	 ),
(	46861	 ),
(	46885	 ),
(	46909	 ),
(	46933	 ),
(	46958	 ),
(	46982	 ),
(	47006	 ),
(	47030	 ),
(	47055	 ),
(	47079	 ),
(	47103	 ),
(	47127	 ),
(	47152	 ),
(	47176	 ),
(	47200	 ),
(	47224	 ),
(	47248	 ),
(	47273	 ),
(	47297	 ),
(	47321	 ),
(	47345	 ),
(	47370	 ),
(	47394	 ),
(	47418	 ),
(	47442	 ),
(	47467	 ),
(	47491	 ),
(	47515	 ),
(	47539	 ),
(	47564	 ),
(	47588	 ),
(	47612	 ),
(	47636	 ),
(	47661	 ),
(	47685	 ),
(	47709	 ),
(	47733	 ),
(	47758	 ),
(	47782	 ),
(	47806	 ),
(	47830	 ),
(	47855	 ),
(	47879	 ),
(	47903	 ),
(	47927	 ),
(	47952	 ),
(	47976	 ),
(	48000	 ),
(	48024	 ),
(	48048	 ),
(	48073	 ),
(	48097	 ),
(	48121	 ),
(	48145	 ),
(	48170	 ),
(	48194	 ),
(	48218	 ),
(	48242	 ),
(	48267	 ),
(	48291	 ),
(	48315	 ),
(	48339	 ),
(	48364	 ),
(	48388	 ),
(	48412	 ),
(	48436	 ),
(	48461	 ),
(	48485	 ),
(	48509	 ),
(	48533	 ),
(	48558	 ),
(	48582	 ),
(	48606	 ),
(	48630	 ),
(	48655	 ),
(	48679	 ),
(	48703	 ),
(	48727	 ),
(	48752	 ),
(	48776	 ),
(	48800	 ),
(	48824	 ),
(	48848	 ),
(	48873	 ),
(	48897	 ),
(	48921	 ),
(	48945	 ),
(	48970	 ),
(	48994	 ),
(	49018	 ),
(	49042	 ),
(	49067	 ),
(	49091	 ),
(	49115	 ),
(	49139	 ),
(	49164	 ),
(	49188	 ),
(	49212	 ),
(	49236	 ),
(	49261	 ),
(	49285	 ),
(	49309	 ),
(	49333	 ),
(	49358	 ),
(	49382	 ),
(	49406	 ),
(	49430	 ),
(	49455	 ),
(	49479	 ),
(	49503	 ),
(	49527	 ),
(	49552	 ),
(	49576	 ),
(	49600	 ),
(	49624	 ),
(	49648	 ),
(	49673	 ),
(	49697	 ),
(	49721	 ),
(	49745	 ),
(	49770	 ),
(	49794	 ),
(	49818	 ),
(	49842	 ),
(	49867	 ),
(	49891	 ),
(	49915	 ),
(	49939	 ),
(	49964	 ),
(	49988	 ),
(	50012	 ),
(	50036	 ),
(	50061	 ),
(	50085	 ),
(	50109	 ),
(	50133	 ),
(	50158	 ),
(	50182	 ),
(	50206	 ),
(	50230	 ),
(	50255	 ),
(	50279	 ),
(	50303	 ),
(	50327	 ),
(	50352	 ),
(	50376	 ),
(	50400	 ),
(	50424	 ),
(	50448	 ),
(	50473	 ),
(	50497	 ),
(	50521	 ),
(	50545	 ),
(	50570	 ),
(	50594	 ),
(	50618	 ),
(	50642	 ),
(	50667	 ),
(	50691	 ),
(	50715	 ),
(	50739	 ),
(	50764	 ),
(	50788	 ),
(	50812	 ),
(	50836	 ),
(	50861	 ),
(	50885	 ),
(	50909	 ),
(	50933	 ),
(	50958	 ),
(	50982	 ),
(	51006	 ),
(	51030	 ),
(	51055	 ),
(	51079	 ),
(	51103	 ),
(	51127	 ),
(	51152	 ),
(	51176	 ),
(	51200	 ),
(	51224	 ),
(	51248	 ),
(	51273	 ),
(	51297	 ),
(	51321	 ),
(	51345	 ),
(	51370	 ),
(	51394	 ),
(	51418	 ),
(	51442	 ),
(	51467	 ),
(	51491	 ),
(	51515	 ),
(	51539	 ),
(	51564	 ),
(	51588	 ),
(	51612	 ),
(	51636	 ),
(	51661	 ),
(	51685	 ),
(	51709	 ),
(	51733	 ),
(	51758	 ),
(	51782	 ),
(	51806	 ),
(	51830	 ),
(	51855	 ),
(	51879	 ),
(	51903	 ),
(	51927	 ),
(	51952	 ),
(	51976	 ),
(	52000	 ),
(	52024	 ),
(	52048	 ),
(	52073	 ),
(	52097	 ),
(	52121	 ),
(	52145	 ),
(	52170	 ),
(	52194	 ),
(	52218	 ),
(	52242	 ),
(	52267	 ),
(	52291	 ),
(	52315	 ),
(	52339	 ),
(	52364	 ),
(	52388	 ),
(	52412	 ),
(	52436	 ),
(	52461	 ),
(	52485	 ),
(	52509	 ),
(	52533	 ),
(	52558	 ),
(	52582	 ),
(	52606	 ),
(	52630	 ),
(	52655	 ),
(	52679	 ),
(	52703	 ),
(	52727	 ),
(	52752	 ),
(	52776	 ),
(	52800	 ),
(	52824	 ),
(	52848	 ),
(	52873	 ),
(	52897	 ),
(	52921	 ),
(	52945	 ),
(	52970	 ),
(	52994	 ),
(	53018	 ),
(	53042	 ),
(	53067	 ),
(	53091	 ),
(	53115	 ),
(	53139	 ),
(	53164	 ),
(	53188	 ),
(	53212	 ),
(	53236	 ),
(	53261	 ),
(	53285	 ),
(	53309	 ),
(	53333	 ),
(	53358	 ),
(	53382	 ),
(	53406	 ),
(	53430	 ),
(	53455	 ),
(	53479	 ),
(	53503	 ),
(	53527	 ),
(	53552	 ),
(	53576	 ),
(	53600	 ),
(	53624	 ),
(	53648	 ),
(	53673	 ),
(	53697	 ),
(	53721	 ),
(	53745	 ),
(	53770	 ),
(	53794	 ),
(	53818	 ),
(	53842	 ),
(	53867	 ),
(	53891	 ),
(	53915	 ),
(	53939	 ),
(	53964	 ),
(	53988	 ),
(	54012	 ),
(	54036	 ),
(	54061	 ),
(	54085	 ),
(	54109	 ),
(	54133	 ),
(	54158	 ),
(	54182	 ),
(	54206	 ),
(	54230	 ),
(	54255	 ),
(	54279	 ),
(	54303	 ),
(	54327	 ),
(	54352	 ),
(	54376	 ),
(	54400	 ),
(	54424	 ),
(	54448	 ),
(	54473	 ),
(	54497	 ),
(	54521	 ),
(	54545	 ),
(	54570	 ),
(	54594	 ),
(	54618	 ),
(	54642	 ),
(	54667	 ),
(	54691	 ),
(	54715	 ),
(	54739	 ),
(	54764	 ),
(	54788	 ),
(	54812	 ),
(	54836	 ),
(	54861	 ),
(	54885	 ),
(	54909	 ),
(	54933	 ),
(	54958	 ),
(	54982	 ),
(	55006	 ),
(	55030	 ),
(	55055	 ),
(	55079	 ),
(	55103	 ),
(	55127	 ),
(	55152	 ),
(	55176	 ),
(	55200	 ),
(	55224	 ),
(	55248	 ),
(	55273	 ),
(	55297	 ),
(	55321	 ),
(	55345	 ),
(	55370	 ),
(	55394	 ),
(	55418	 ),
(	55442	 ),
(	55467	 ),
(	55491	 ),
(	55515	 ),
(	55539	 ),
(	55564	 ),
(	55588	 ),
(	55612	 ),
(	55636	 ),
(	55661	 ),
(	55685	 ),
(	55709	 ),
(	55733	 ),
(	55758	 ),
(	55782	 ),
(	55806	 ),
(	55830	 ),
(	55855	 ),
(	55879	 ),
(	55903	 ),
(	55927	 ),
(	55952	 ),
(	55976	 ),
(	56000	 ),
(	56024	 ),
(	56048	 ),
(	56073	 ),
(	56097	 ),
(	56121	 ),
(	56145	 ),
(	56170	 ),
(	56194	 ),
(	56218	 ),
(	56242	 ),
(	56267	 ),
(	56291	 ),
(	56315	 ),
(	56339	 ),
(	56364	 ),
(	56388	 ),
(	56412	 ),
(	56436	 ),
(	56461	 ),
(	56485	 ),
(	56509	 ),
(	56533	 ),
(	56558	 ),
(	56582	 ),
(	56606	 ),
(	56630	 ),
(	56655	 ),
(	56679	 ),
(	56703	 ),
(	56727	 ),
(	56752	 ),
(	56776	 ),
(	56800	 ),
(	56824	 ),
(	56848	 ),
(	56873	 ),
(	56897	 ),
(	56921	 ),
(	56945	 ),
(	56970	 ),
(	56994	 ),
(	57018	 ),
(	57042	 ),
(	57067	 ),
(	57091	 ),
(	57115	 ),
(	57139	 ),
(	57164	 ),
(	57188	 ),
(	57212	 ),
(	57236	 ),
(	57261	 ),
(	57285	 ),
(	57309	 ),
(	57333	 ),
(	57358	 ),
(	57382	 ),
(	57406	 ),
(	57430	 ),
(	57455	 ),
(	57479	 ),
(	57503	 ),
(	57527	 ),
(	57552	 ),
(	57576	 ),
(	57600	 ),
(	57624	 ),
(	57648	 ),
(	57673	 ),
(	57697	 ),
(	57721	 ),
(	57745	 ),
(	57770	 ),
(	57794	 ),
(	57818	 ),
(	57842	 ),
(	57867	 ),
(	57891	 ),
(	57915	 ),
(	57939	 ),
(	57964	 ),
(	57988	 ),
(	58012	 ),
(	58036	 ),
(	58061	 ),
(	58085	 ),
(	58109	 ),
(	58133	 ),
(	58158	 ),
(	58182	 ),
(	58206	 ),
(	58230	 ),
(	58255	 ),
(	58279	 ),
(	58303	 ),
(	58327	 ),
(	58352	 ),
(	58376	 ),
(	58400	 ),
(	58424	 ),
(	58448	 ),
(	58473	 ),
(	58497	 ),
(	58521	 ),
(	58545	 ),
(	58570	 ),
(	58594	 ),
(	58618	 ),
(	58642	 ),
(	58667	 ),
(	58691	 ),
(	58715	 ),
(	58739	 ),
(	58764	 ),
(	58788	 ),
(	58812	 ),
(	58836	 ),
(	58861	 ),
(	58885	 ),
(	58909	 ),
(	58933	 ),
(	58958	 ),
(	58982	 ),
(	59006	 ),
(	59030	 ),
(	59055	 ),
(	59079	 ),
(	59103	 ),
(	59127	 ),
(	59152	 ),
(	59176	 ),
(	59200	 ),
(	59224	 ),
(	59248	 ),
(	59273	 ),
(	59297	 ),
(	59321	 ),
(	59345	 ),
(	59370	 ),
(	59394	 ),
(	59418	 ),
(	59442	 ),
(	59467	 ),
(	59491	 ),
(	59515	 ),
(	59539	 ),
(	59564	 ),
(	59588	 ),
(	59612	 ),
(	59636	 ),
(	59661	 ),
(	59685	 ),
(	59709	 ),
(	59733	 ),
(	59758	 ),
(	59782	 ),
(	59806	 ),
(	59830	 ),
(	59855	 ),
(	59879	 ),
(	59903	 ),
(	59927	 ),
(	59952	 ),
(	59976	 ),
(	60000	 ),
(	60024	 ),
(	60048	 ),
(	60073	 ),
(	60097	 ),
(	60121	 ),
(	60145	 ),
(	60170	 ),
(	60194	 ),
(	60218	 ),
(	60242	 ),
(	60267	 ),
(	60291	 ),
(	60315	 ),
(	60339	 ),
(	60364	 ),
(	60388	 ),
(	60412	 ),
(	60436	 ),
(	60461	 ),
(	60485	 ),
(	60509	 ),
(	60533	 ),
(	60558	 ),
(	60582	 ),
(	60606	 ),
(	60630	 ),
(	60655	 ),
(	60679	 ),
(	60703	 ),
(	60727	 ),
(	60752	 ),
(	60776	 ),
(	60800	 ),
(	60824	 ),
(	60848	 ),
(	60873	 ),
(	60897	 ),
(	60921	 ),
(	60945	 ),
(	60970	 ),
(	60994	 ),
(	61018	 ),
(	61042	 ),
(	61067	 ),
(	61091	 ),
(	61115	 ),
(	61139	 ),
(	61164	 ),
(	61188	 ),
(	61212	 ),
(	61236	 ),
(	61261	 ),
(	61285	 ),
(	61309	 ),
(	61333	 ),
(	61358	 ),
(	61382	 ),
(	61406	 ),
(	61430	 ),
(	61455	 ),
(	61479	 ),
(	61503	 ),
(	61527	 ),
(	61552	 ),
(	61576	 ),
(	61600	 ),
(	61624	 ),
(	61648	 ),
(	61673	 ),
(	61697	 ),
(	61721	 ),
(	61745	 ),
(	61770	 ),
(	61794	 ),
(	61818	 ),
(	61842	 ),
(	61867	 ),
(	61891	 ),
(	61915	 ),
(	61939	 ),
(	61964	 ),
(	61988	 ),
(	62012	 ),
(	62036	 ),
(	62061	 ),
(	62085	 ),
(	62109	 ),
(	62133	 ),
(	62158	 ),
(	62182	 ),
(	62206	 ),
(	62230	 ),
(	62255	 ),
(	62279	 ),
(	62303	 ),
(	62327	 ),
(	62352	 ),
(	62376	 ),
(	62400	 ),
(	62424	 ),
(	62448	 ),
(	62473	 ),
(	62497	 ),
(	62521	 ),
(	62545	 ),
(	62570	 ),
(	62594	 ),
(	62618	 ),
(	62642	 ),
(	62667	 ),
(	62691	 ),
(	62715	 ),
(	62739	 ),
(	62764	 ),
(	62788	 ),
(	62812	 ),
(	62836	 ),
(	62861	 ),
(	62885	 ),
(	62909	 ),
(	62933	 ),
(	62958	 ),
(	62982	 ),
(	63006	 ),
(	63030	 ),
(	63055	 ),
(	63079	 ),
(	63103	 ),
(	63127	 ),
(	63152	 ),
(	63176	 ),
(	63200	 ),
(	63224	 ),
(	63248	 ),
(	63273	 ),
(	63297	 ),
(	63321	 ),
(	63345	 ),
(	63370	 ),
(	63394	 ),
(	63418	 ),
(	63442	 ),
(	63467	 ),
(	63491	 ),
(	63515	 ),
(	63539	 ),
(	63564	 ),
(	63588	 ),
(	63612	 ),
(	63636	 ),
(	63661	 ),
(	63685	 ),
(	63709	 ),
(	63733	 ),
(	63758	 ),
(	63782	 ),
(	63806	 ),
(	63830	 ),
(	63855	 ),
(	63879	 ),
(	63903	 ),
(	63927	 ),
(	63952	 ),
(	63976	 ),
(	64000	 ),
(	64024	 ),
(	64048	 ),
(	64073	 ),
(	64097	 ),
(	64121	 ),
(	64145	 ),
(	64170	 ),
(	64194	 ),
(	64218	 ),
(	64242	 ),
(	64267	 ),
(	64291	 ),
(	64315	 ),
(	64339	 ),
(	64364	 ),
(	64388	 ),
(	64412	 ),
(	64436	 ),
(	64461	 ),
(	64485	 ),
(	64509	 ),
(	64533	 ),
(	64558	 ),
(	64582	 ),
(	64606	 ),
(	64630	 ),
(	64655	 ),
(	64679	 ),
(	64703	 ),
(	64727	 ),
(	64752	 ),
(	64776	 ),
(	64800	 ),
(	64824	 ),
(	64848	 ),
(	64873	 ),
(	64897	 ),
(	64921	 ),
(	64945	 ),
(	64970	 ),
(	64994	 ),
(	65018	 ),
(	65042	 ),
(	65067	 ),
(	65091	 ),
(	65115	 ),
(	65139	 ),
(	65164	 ),
(	65188	 ),
(	65212	 ),
(	65236	 ),
(	65261	 ),
(	65285	 ),
(	65309	 ),
(	65333	 ),
(	65358	 ),
(	65382	 ),
(	65406	 ),
(	65430	 ),
(	65455	 ),
(	65479	 ),
(	65503	 ),
(	65527	 ),
(	65552	 ),
(	65576	 ),
(	65600	 ),
(	65624	 ),
(	65648	 ),
(	65673	 ),
(	65697	 ),
(	65721	 ),
(	65745	 ),
(	65770	 ),
(	65794	 ),
(	65818	 ),
(	65842	 ),
(	65867	 ),
(	65891	 ),
(	65915	 ),
(	65939	 ),
(	65964	 ),
(	65988	 ),
(	66012	 ),
(	66036	 ),
(	66061	 ),
(	66085	 ),
(	66109	 ),
(	66133	 ),
(	66158	 ),
(	66182	 ),
(	66206	 ),
(	66230	 ),
(	66255	 ),
(	66279	 ),
(	66303	 ),
(	66327	 ),
(	66352	 ),
(	66376	 ),
(	66400	 ),
(	66424	 ),
(	66448	 ),
(	66473	 ),
(	66497	 ),
(	66521	 ),
(	66545	 ),
(	66570	 ),
(	66594	 ),
(	66618	 ),
(	66642	 ),
(	66667	 ),
(	66691	 ),
(	66715	 ),
(	66739	 ),
(	66764	 ),
(	66788	 ),
(	66812	 ),
(	66836	 ),
(	66861	 ),
(	66885	 ),
(	66909	 ),
(	66933	 ),
(	66958	 ),
(	66982	 ),
(	67006	 ),
(	67030	 ),
(	67055	 ),
(	67079	 ),
(	67103	 ),
(	67127	 ),
(	67152	 ),
(	67176	 ),
(	67200	 ),
(	67224	 ),
(	67248	 ),
(	67273	 ),
(	67297	 ),
(	67321	 ),
(	67345	 ),
(	67370	 ),
(	67394	 ),
(	67418	 ),
(	67442	 ),
(	67467	 ),
(	67491	 ),
(	67515	 ),
(	67539	 ),
(	67564	 ),
(	67588	 ),
(	67612	 ),
(	67636	 ),
(	67661	 ),
(	67685	 ),
(	67709	 ),
(	67733	 ),
(	67758	 ),
(	67782	 ),
(	67806	 ),
(	67830	 ),
(	67855	 ),
(	67879	 ),
(	67903	 ),
(	67927	 ),
(	67952	 ),
(	67976	 ),
(	68000	 ),
(	68024	 ),
(	68048	 ),
(	68073	 ),
(	68097	 ),
(	68121	 ),
(	68145	 ),
(	68170	 ),
(	68194	 ),
(	68218	 ),
(	68242	 ),
(	68267	 ),
(	68291	 ),
(	68315	 ),
(	68339	 ),
(	68364	 ),
(	68388	 ),
(	68412	 ),
(	68436	 ),
(	68461	 ),
(	68485	 ),
(	68509	 ),
(	68533	 ),
(	68558	 ),
(	68582	 ),
(	68606	 ),
(	68630	 ),
(	68655	 ),
(	68679	 ),
(	68703	 ),
(	68727	 ),
(	68752	 ),
(	68776	 ),
(	68800	 ),
(	68824	 ),
(	68848	 ),
(	68873	 ),
(	68897	 ),
(	68921	 ),
(	68945	 ),
(	68970	 ),
(	68994	 ),
(	69018	 ),
(	69042	 ),
(	69067	 ),
(	69091	 ),
(	69115	 ),
(	69139	 ),
(	69164	 ),
(	69188	 ),
(	69212	 ),
(	69236	 ),
(	69261	 ),
(	69285	 ),
(	69309	 ),
(	69333	 ),
(	69358	 ),
(	69382	 ),
(	69406	 ),
(	69430	 ),
(	69455	 ),
(	69479	 ),
(	69503	 ),
(	69527	 ),
(	69552	 ),
(	69576	 ),
(	69600	 ),
(	69624	 ),
(	69648	 ),
(	69673	 ),
(	69697	 ),
(	69721	 ),
(	69745	 ),
(	69770	 ),
(	69794	 ),
(	69818	 ),
(	69842	 ),
(	69867	 ),
(	69891	 ),
(	69915	 ),
(	69939	 ),
(	69964	 ),
(	69988	 ),
(	70012	 ),
(	70036	 ),
(	70061	 ),
(	70085	 ),
(	70109	 ),
(	70133	 ),
(	70158	 ),
(	70182	 ),
(	70206	 ),
(	70230	 ),
(	70255	 ),
(	70279	 ),
(	70303	 ),
(	70327	 ),
(	70352	 ),
(	70376	 ),
(	70400	 ),
(	70424	 ),
(	70448	 ),
(	70473	 ),
(	70497	 ),
(	70521	 ),
(	70545	 ),
(	70570	 ),
(	70594	 ),
(	70618	 ),
(	70642	 ),
(	70667	 ),
(	70691	 ),
(	70715	 ),
(	70739	 ),
(	70764	 ),
(	70788	 ),
(	70812	 ),
(	70836	 ),
(	70861	 ),
(	70885	 ),
(	70909	 ),
(	70933	 ),
(	70958	 ),
(	70982	 ),
(	71006	 ),
(	71030	 ),
(	71055	 ),
(	71079	 ),
(	71103	 ),
(	71127	 ),
(	71152	 ),
(	71176	 ),
(	71200	 ),
(	71224	 ),
(	71248	 ),
(	71273	 ),
(	71297	 ),
(	71321	 ),
(	71345	 ),
(	71370	 ),
(	71394	 ),
(	71418	 ),
(	71442	 ),
(	71467	 ),
(	71491	 ),
(	71515	 ),
(	71539	 ),
(	71564	 ),
(	71588	 ),
(	71612	 ),
(	71636	 ),
(	71661	 ),
(	71685	 ),
(	71709	 ),
(	71733	 ),
(	71758	 ),
(	71782	 ),
(	71806	 ),
(	71830	 ),
(	71855	 ),
(	71879	 ),
(	71903	 ),
(	71927	 ),
(	71952	 ),
(	71976	 ),
(	72000	 ),
(	72024	 ),
(	72048	 ),
(	72073	 ),
(	72097	 ),
(	72121	 ),
(	72145	 ),
(	72170	 ),
(	72194	 ),
(	72218	 ),
(	72242	 ),
(	72267	 ),
(	72291	 ),
(	72315	 ),
(	72339	 ),
(	72364	 ),
(	72388	 ),
(	72412	 ),
(	72436	 ),
(	72461	 ),
(	72485	 ),
(	72509	 ),
(	72533	 ),
(	72558	 ),
(	72582	 ),
(	72606	 ),
(	72630	 ),
(	72655	 ),
(	72679	 ),
(	72703	 ),
(	72727	 ),
(	72752	 ),
(	72776	 ),
(	72800	 ),
(	72824	 ),
(	72848	 ),
(	72873	 ),
(	72897	 ),
(	72921	 ),
(	72945	 ),
(	72970	 ),
(	72994	 ),
(	73018	 ),
(	73042	 ),
(	73067	 ),
(	73091	 ),
(	73115	 ),
(	73139	 ),
(	73164	 ),
(	73188	 ),
(	73212	 ),
(	73236	 ),
(	73261	 ),
(	73285	 ),
(	73309	 ),
(	73333	 ),
(	73358	 ),
(	73382	 ),
(	73406	 ),
(	73430	 ),
(	73455	 ),
(	73479	 ),
(	73503	 ),
(	73527	 ),
(	73552	 ),
(	73576	 ),
(	73600	 ),
(	73624	 ),
(	73648	 ),
(	73673	 ),
(	73697	 ),
(	73721	 ),
(	73745	 ),
(	73770	 ),
(	73794	 ),
(	73818	 ),
(	73842	 ),
(	73867	 ),
(	73891	 ),
(	73915	 ),
(	73939	 ),
(	73964	 ),
(	73988	 ),
(	74012	 ),
(	74036	 ),
(	74061	 ),
(	74085	 ),
(	74109	 ),
(	74133	 ),
(	74158	 ),
(	74182	 ),
(	74206	 ),
(	74230	 ),
(	74255	 ),
(	74279	 ),
(	74303	 ),
(	74327	 ),
(	74352	 ),
(	74376	 ),
(	74400	 ),
(	74424	 ),
(	74448	 ),
(	74473	 ),
(	74497	 ),
(	74521	 ),
(	74545	 ),
(	74570	 ),
(	74594	 ),
(	74618	 ),
(	74642	 ),
(	74667	 ),
(	74691	 ),
(	74715	 ),
(	74739	 ),
(	74764	 ),
(	74788	 ),
(	74812	 ),
(	74836	 ),
(	74861	 ),
(	74885	 ),
(	74909	 ),
(	74933	 ),
(	74958	 ),
(	74982	 ),
(	75006	 ),
(	75030	 ),
(	75055	 ),
(	75079	 ),
(	75103	 ),
(	75127	 ),
(	75152	 ),
(	75176	 ),
(	75200	 ),
(	75224	 ),
(	75248	 ),
(	75273	 ),
(	75297	 ),
(	75321	 ),
(	75345	 ),
(	75370	 ),
(	75394	 ),
(	75418	 ),
(	75442	 ),
(	75467	 ),
(	75491	 ),
(	75515	 ),
(	75539	 ),
(	75564	 ),
(	75588	 ),
(	75612	 ),
(	75636	 ),
(	75661	 ),
(	75685	 ),
(	75709	 ),
(	75733	 ),
(	75758	 ),
(	75782	 ),
(	75806	 ),
(	75830	 ),
(	75855	 ),
(	75879	 ),
(	75903	 ),
(	75927	 ),
(	75952	 ),
(	75976	 ),
(	76000	 ),
(	76024	 ),
(	76048	 ),
(	76073	 ),
(	76097	 ),
(	76121	 ),
(	76145	 ),
(	76170	 ),
(	76194	 ),
(	76218	 ),
(	76242	 ),
(	76267	 ),
(	76291	 ),
(	76315	 ),
(	76339	 ),
(	76364	 ),
(	76388	 ),
(	76412	 ),
(	76436	 ),
(	76461	 ),
(	76485	 ),
(	76509	 ),
(	76533	 ),
(	76558	 ),
(	76582	 ),
(	76606	 ),
(	76630	 ),
(	76655	 ),
(	76679	 ),
(	76703	 ),
(	76727	 ),
(	76752	 ),
(	76776	 ),
(	76800	 ),
(	76824	 ),
(	76848	 ),
(	76873	 ),
(	76897	 ),
(	76921	 ),
(	76945	 ),
(	76970	 ),
(	76994	 ),
(	77018	 ),
(	77042	 ),
(	77067	 ),
(	77091	 ),
(	77115	 ),
(	77139	 ),
(	77164	 ),
(	77188	 ),
(	77212	 ),
(	77236	 ),
(	77261	 ),
(	77285	 ),
(	77309	 ),
(	77333	 ),
(	77358	 ),
(	77382	 ),
(	77406	 ),
(	77430	 ),
(	77455	 ),
(	77479	 ),
(	77503	 ),
(	77527	 ),
(	77552	 ),
(	77576	 ),
(	77600	 ),
(	77624	 ),
(	77648	 ),
(	77673	 ),
(	77697	 ),
(	77721	 ),
(	77745	 ),
(	77770	 ),
(	77794	 ),
(	77818	 ),
(	77842	 ),
(	77867	 ),
(	77891	 ),
(	77915	 ),
(	77939	 ),
(	77964	 ),
(	77988	 ),
(	78012	 ),
(	78036	 ),
(	78061	 ),
(	78085	 ),
(	78109	 ),
(	78133	 ),
(	78158	 ),
(	78182	 ),
(	78206	 ),
(	78230	 ),
(	78255	 ),
(	78279	 ),
(	78303	 ),
(	78327	 ),
(	78352	 ),
(	78376	 ),
(	78400	 ),
(	78424	 ),
(	78448	 ),
(	78473	 ),
(	78497	 ),
(	78521	 ),
(	78545	 ),
(	78570	 ),
(	78594	 ),
(	78618	 ),
(	78642	 ),
(	78667	 ),
(	78691	 ),
(	78715	 ),
(	78739	 ),
(	78764	 ),
(	78788	 ),
(	78812	 ),
(	78836	 ),
(	78861	 ),
(	78885	 ),
(	78909	 ),
(	78933	 ),
(	78958	 ),
(	78982	 ),
(	79006	 ),
(	79030	 ),
(	79055	 ),
(	79079	 ),
(	79103	 ),
(	79127	 ),
(	79152	 ),
(	79176	 ),
(	79200	 ),
(	79224	 ),
(	79248	 ),
(	79273	 ),
(	79297	 ),
(	79321	 ),
(	79345	 ),
(	79370	 ),
(	79394	 ),
(	79418	 ),
(	79442	 ),
(	79467	 ),
(	79491	 ),
(	79515	 ),
(	79539	 ),
(	79564	 ),
(	79588	 ),
(	79612	 ),
(	79636	 ),
(	79661	 ),
(	79685	 ),
(	79709	 ),
(	79733	 ),
(	79758	 ),
(	79782	 ),
(	79806	 ),
(	79830	 ),
(	79855	 ),
(	79879	 ),
(	79903	 ),
(	79927	 ),
(	79952	 ),
(	79976	 ),
(	80000	 ),
(	80024	 ),
(	80048	 ),
(	80073	 ),
(	80097	 ),
(	80121	 ),
(	80145	 ),
(	80170	 ),
(	80194	 ),
(	80218	 ),
(	80242	 ),
(	80267	 ),
(	80291	 ),
(	80315	 ),
(	80339	 ),
(	80364	 ),
(	80388	 ),
(	80412	 ),
(	80436	 ),
(	80461	 ),
(	80485	 ),
(	80509	 ),
(	80533	 ),
(	80558	 ),
(	80582	 ),
(	80606	 ),
(	80630	 ),
(	80655	 ),
(	80679	 ),
(	80703	 ),
(	80727	 ),
(	80752	 ),
(	80776	 ),
(	80800	 ),
(	80824	 ),
(	80848	 ),
(	80873	 ),
(	80897	 ),
(	80921	 ),
(	80945	 ),
(	80970	 ),
(	80994	 ),
(	81018	 ),
(	81042	 ),
(	81067	 ),
(	81091	 ),
(	81115	 ),
(	81139	 ),
(	81164	 ),
(	81188	 ),
(	81212	 ),
(	81236	 ),
(	81261	 ),
(	81285	 ),
(	81309	 ),
(	81333	 ),
(	81358	 ),
(	81382	 ),
(	81406	 ),
(	81430	 ),
(	81455	 ),
(	81479	 ),
(	81503	 ),
(	81527	 ),
(	81552	 ),
(	81576	 ),
(	81600	 ),
(	81624	 ),
(	81648	 ),
(	81673	 ),
(	81697	 ),
(	81721	 ),
(	81745	 ),
(	81770	 ),
(	81794	 ),
(	81818	 ),
(	81842	 ),
(	81867	 ),
(	81891	 ),
(	81915	 ),
(	81939	 ),
(	81964	 ),
(	81988	 ),
(	82012	 ),
(	82036	 ),
(	82061	 ),
(	82085	 ),
(	82109	 ),
(	82133	 ),
(	82158	 ),
(	82182	 ),
(	82206	 ),
(	82230	 ),
(	82255	 ),
(	82279	 ),
(	82303	 ),
(	82327	 ),
(	82352	 ),
(	82376	 ),
(	82400	 ),
(	82424	 ),
(	82448	 ),
(	82473	 ),
(	82497	 ),
(	82521	 ),
(	82545	 ),
(	82570	 ),
(	82594	 ),
(	82618	 ),
(	82642	 ),
(	82667	 ),
(	82691	 ),
(	82715	 ),
(	82739	 ),
(	82764	 ),
(	82788	 ),
(	82812	 ),
(	82836	 ),
(	82861	 ),
(	82885	 ),
(	82909	 ),
(	82933	 ),
(	82958	 ),
(	82982	 ),
(	83006	 ),
(	83030	 ),
(	83055	 ),
(	83079	 ),
(	83103	 ),
(	83127	 ),
(	83152	 ),
(	83176	 ),
(	83200	 ),
(	83224	 ),
(	83248	 ),
(	83273	 ),
(	83297	 ),
(	83321	 ),
(	83345	 ),
(	83370	 ),
(	83394	 ),
(	83418	 ),
(	83442	 ),
(	83467	 ),
(	83491	 ),
(	83515	 ),
(	83539	 ),
(	83564	 ),
(	83588	 ),
(	83612	 ),
(	83636	 ),
(	83661	 ),
(	83685	 ),
(	83709	 ),
(	83733	 ),
(	83758	 ),
(	83782	 ),
(	83806	 ),
(	83830	 ),
(	83855	 ),
(	83879	 ),
(	83903	 ),
(	83927	 ),
(	83952	 ),
(	83976	 ),
(	84000	 ),
(	84024	 ),
(	84048	 ),
(	84073	 ),
(	84097	 ),
(	84121	 ),
(	84145	 ),
(	84170	 ),
(	84194	 ),
(	84218	 ),
(	84242	 ),
(	84267	 ),
(	84291	 ),
(	84315	 ),
(	84339	 ),
(	84364	 ),
(	84388	 ),
(	84412	 ),
(	84436	 ),
(	84461	 ),
(	84485	 ),
(	84509	 ),
(	84533	 ),
(	84558	 ),
(	84582	 ),
(	84606	 ),
(	84630	 ),
(	84655	 ),
(	84679	 ),
(	84703	 ),
(	84727	 ),
(	84752	 ),
(	84776	 ),
(	84800	 ),
(	84824	 ),
(	84848	 ),
(	84873	 ),
(	84897	 ),
(	84921	 ),
(	84945	 ),
(	84970	 ),
(	84994	 ),
(	85018	 ),
(	85042	 ),
(	85067	 ),
(	85091	 ),
(	85115	 ),
(	85139	 ),
(	85164	 ),
(	85188	 ),
(	85212	 ),
(	85236	 ),
(	85261	 ),
(	85285	 ),
(	85309	 ),
(	85333	 ),
(	85358	 ),
(	85382	 ),
(	85406	 ),
(	85430	 ),
(	85455	 ),
(	85479	 ),
(	85503	 ),
(	85527	 ),
(	85552	 ),
(	85576	 ),
(	85600	 ),
(	85624	 ),
(	85648	 ),
(	85673	 ),
(	85697	 ),
(	85721	 ),
(	85745	 ),
(	85770	 ),
(	85794	 ),
(	85818	 ),
(	85842	 ),
(	85867	 ),
(	85891	 ),
(	85915	 ),
(	85939	 ),
(	85964	 ),
(	85988	 ),
(	86012	 ),
(	86036	 ),
(	86061	 ),
(	86085	 ),
(	86109	 ),
(	86133	 ),
(	86158	 ),
(	86182	 ),
(	86206	 ),
(	86230	 ),
(	86255	 ),
(	86279	 ),
(	86303	 ),
(	86327	 ),
(	86352	 ),
(	86376	 ),
(	86400	 ),
(	86424	 ),
(	86448	 ),
(	86473	 ),
(	86497	 ),
(	86521	 ),
(	86545	 ),
(	86570	 ),
(	86594	 ),
(	86618	 ),
(	86642	 ),
(	86667	 ),
(	86691	 ),
(	86715	 ),
(	86739	 ),
(	86764	 ),
(	86788	 ),
(	86812	 ),
(	86836	 ),
(	86861	 ),
(	86885	 ),
(	86909	 ),
(	86933	 ),
(	86958	 ),
(	86982	 ),
(	87006	 ),
(	87030	 ),
(	87055	 ),
(	87079	 ),
(	87103	 ),
(	87127	 ),
(	87152	 ),
(	87176	 ),
(	87200	 ),
(	87224	 ),
(	87248	 ),
(	87273	 ),
(	87297	 ),
(	87321	 ),
(	87345	 ),
(	87370	 ),
(	87394	 ),
(	87418	 ),
(	87442	 ),
(	87467	 ),
(	87491	 ),
(	87515	 ),
(	87539	 ),
(	87564	 ),
(	87588	 ),
(	87612	 ),
(	87636	 ),
(	87661	 ),
(	87685	 ),
(	87709	 ),
(	87733	 ),
(	87758	 ),
(	87782	 ),
(	87806	 ),
(	87830	 ),
(	87855	 ),
(	87879	 ),
(	87903	 ),
(	87927	 ),
(	87952	 ),
(	87976	 ),
(	88000	 ),
(	88024	 ),
(	88048	 ),
(	88073	 ),
(	88097	 ),
(	88121	 ),
(	88145	 ),
(	88170	 ),
(	88194	 ),
(	88218	 ),
(	88242	 ),
(	88267	 ),
(	88291	 ),
(	88315	 ),
(	88339	 ),
(	88364	 ),
(	88388	 ),
(	88412	 ),
(	88436	 ),
(	88461	 ),
(	88485	 ),
(	88509	 ),
(	88533	 ),
(	88558	 ),
(	88582	 ),
(	88606	 ),
(	88630	 ),
(	88655	 ),
(	88679	 ),
(	88703	 ),
(	88727	 ),
(	88752	 ),
(	88776	 ),
(	88800	 ),
(	88824	 ),
(	88848	 ),
(	88873	 ),
(	88897	 ),
(	88921	 ),
(	88945	 ),
(	88970	 ),
(	88994	 ),
(	89018	 ),
(	89042	 ),
(	89067	 ),
(	89091	 ),
(	89115	 ),
(	89139	 ),
(	89164	 ),
(	89188	 ),
(	89212	 ),
(	89236	 ),
(	89261	 ),
(	89285	 ),
(	89309	 ),
(	89333	 ),
(	89358	 ),
(	89382	 ),
(	89406	 ),
(	89430	 ),
(	89455	 ),
(	89479	 ),
(	89503	 ),
(	89527	 ),
(	89552	 ),
(	89576	 ),
(	89600	 ),
(	89624	 ),
(	89648	 ),
(	89673	 ),
(	89697	 ),
(	89721	 ),
(	89745	 ),
(	89770	 ),
(	89794	 ),
(	89818	 ),
(	89842	 ),
(	89867	 ),
(	89891	 ),
(	89915	 ),
(	89939	 ),
(	89964	 ),
(	89988	 ),
(	90012	 ),
(	90036	 ),
(	90061	 ),
(	90085	 ),
(	90109	 ),
(	90133	 ),
(	90158	 ),
(	90182	 ),
(	90206	 ),
(	90230	 ),
(	90255	 ),
(	90279	 ),
(	90303	 ),
(	90327	 ),
(	90352	 ),
(	90376	 ),
(	90400	 ),
(	90424	 ),
(	90448	 ),
(	90473	 ),
(	90497	 ),
(	90521	 ),
(	90545	 ),
(	90570	 ),
(	90594	 ),
(	90618	 ),
(	90642	 ),
(	90667	 ),
(	90691	 ),
(	90715	 ),
(	90739	 ),
(	90764	 ),
(	90788	 ),
(	90812	 ),
(	90836	 ),
(	90861	 ),
(	90885	 ),
(	90909	 ),
(	90933	 ),
(	90958	 ),
(	90982	 ),
(	91006	 ),
(	91030	 ),
(	91055	 ),
(	91079	 ),
(	91103	 ),
(	91127	 ),
(	91152	 ),
(	91176	 ),
(	91200	 ),
(	91224	 ),
(	91248	 ),
(	91273	 ),
(	91297	 ),
(	91321	 ),
(	91345	 ),
(	91370	 ),
(	91394	 ),
(	91418	 ),
(	91442	 ),
(	91467	 ),
(	91491	 ),
(	91515	 ),
(	91539	 ),
(	91564	 ),
(	91588	 ),
(	91612	 ),
(	91636	 ),
(	91661	 ),
(	91685	 ),
(	91709	 ),
(	91733	 ),
(	91758	 ),
(	91782	 ),
(	91806	 ),
(	91830	 ),
(	91855	 ),
(	91879	 ),
(	91903	 ),
(	91927	 ),
(	91952	 ),
(	91976	 ),
(	92000	 ),
(	92024	 ),
(	92048	 ),
(	92073	 ),
(	92097	 ),
(	92121	 ),
(	92145	 ),
(	92170	 ),
(	92194	 ),
(	92218	 ),
(	92242	 ),
(	92267	 ),
(	92291	 ),
(	92315	 ),
(	92339	 ),
(	92364	 ),
(	92388	 ),
(	92412	 ),
(	92436	 ),
(	92461	 ),
(	92485	 ),
(	92509	 ),
(	92533	 ),
(	92558	 ),
(	92582	 ),
(	92606	 ),
(	92630	 ),
(	92655	 ),
(	92679	 ),
(	92703	 ),
(	92727	 ),
(	92752	 ),
(	92776	 ),
(	92800	 ),
(	92824	 ),
(	92848	 ),
(	92873	 ),
(	92897	 ),
(	92921	 ),
(	92945	 ),
(	92970	 ),
(	92994	 ),
(	93018	 ),
(	93042	 ),
(	93067	 ),
(	93091	 ),
(	93115	 ),
(	93139	 ),
(	93164	 ),
(	93188	 ),
(	93212	 ),
(	93236	 ),
(	93261	 ),
(	93285	 ),
(	93309	 ),
(	93333	 ),
(	93358	 ),
(	93382	 ),
(	93406	 ),
(	93430	 ),
(	93455	 ),
(	93479	 ),
(	93503	 ),
(	93527	 ),
(	93552	 ),
(	93576	 ),
(	93600	 ),
(	93624	 ),
(	93648	 ),
(	93673	 ),
(	93697	 ),
(	93721	 ),
(	93745	 ),
(	93770	 ),
(	93794	 ),
(	93818	 ),
(	93842	 ),
(	93867	 ),
(	93891	 ),
(	93915	 ),
(	93939	 ),
(	93964	 ),
(	93988	 ),
(	94012	 ),
(	94036	 ),
(	94061	 ),
(	94085	 ),
(	94109	 ),
(	94133	 ),
(	94158	 ),
(	94182	 ),
(	94206	 ),
(	94230	 ),
(	94255	 ),
(	94279	 ),
(	94303	 ),
(	94327	 ),
(	94352	 ),
(	94376	 ),
(	94400	 ),
(	94424	 ),
(	94448	 ),
(	94473	 ),
(	94497	 ),
(	94521	 ),
(	94545	 ),
(	94570	 ),
(	94594	 ),
(	94618	 ),
(	94642	 ),
(	94667	 ),
(	94691	 ),
(	94715	 ),
(	94739	 ),
(	94764	 ),
(	94788	 ),
(	94812	 ),
(	94836	 ),
(	94861	 ),
(	94885	 ),
(	94909	 ),
(	94933	 ),
(	94958	 ),
(	94982	 ),
(	95006	 ),
(	95030	 ),
(	95055	 ),
(	95079	 ),
(	95103	 ),
(	95127	 ),
(	95152	 ),
(	95176	 ),
(	95200	 ),
(	95224	 ),
(	95248	 ),
(	95273	 ),
(	95297	 ),
(	95321	 ),
(	95345	 ),
(	95370	 ),
(	95394	 ),
(	95418	 ),
(	95442	 ),
(	95467	 ),
(	95491	 ),
(	95515	 ),
(	95539	 ),
(	95564	 ),
(	95588	 ),
(	95612	 ),
(	95636	 ),
(	95661	 ),
(	95685	 ),
(	95709	 ),
(	95733	 ),
(	95758	 ),
(	95782	 ),
(	95806	 ),
(	95830	 ),
(	95855	 ),
(	95879	 ),
(	95903	 ),
(	95927	 ),
(	95952	 ),
(	95976	 ),
(	96000	 ),
(	96024	 ),
(	96048	 ),
(	96073	 ),
(	96097	 ),
(	96121	 ),
(	96145	 ),
(	96170	 ),
(	96194	 ),
(	96218	 ),
(	96242	 ),
(	96267	 ),
(	96291	 ),
(	96315	 ),
(	96339	 ),
(	96364	 ),
(	96388	 ),
(	96412	 ),
(	96436	 ),
(	96461	 ),
(	96485	 ),
(	96509	 ),
(	96533	 ),
(	96558	 ),
(	96582	 ),
(	96606	 ),
(	96630	 ),
(	96655	 ),
(	96679	 ),
(	96703	 ),
(	96727	 ),
(	96752	 ),
(	96776	 ),
(	96800	 ),
(	96824	 ),
(	96848	 ),
(	96873	 ),
(	96897	 ),
(	96921	 ),
(	96945	 ),
(	96970	 ),
(	96994	 ),
(	97018	 ),
(	97042	 ),
(	97067	 ),
(	97091	 ),
(	97115	 ),
(	97139	 ),
(	97164	 ),
(	97188	 ),
(	97212	 ),
(	97236	 ),
(	97261	 ),
(	97285	 ),
(	97309	 ),
(	97333	 ),
(	97358	 ),
(	97382	 ),
(	97406	 ),
(	97430	 ),
(	97455	 ),
(	97479	 ),
(	97503	 ),
(	97527	 ),
(	97552	 ),
(	97576	 ),
(	97600	 ),
(	97624	 ),
(	97648	 ),
(	97673	 ),
(	97697	 ),
(	97721	 ),
(	97745	 ),
(	97770	 ),
(	97794	 ),
(	97818	 ),
(	97842	 ),
(	97867	 ),
(	97891	 ),
(	97915	 ),
(	97939	 ),
(	97964	 ),
(	97988	 ),
(	98012	 ),
(	98036	 ),
(	98061	 ),
(	98085	 ),
(	98109	 ),
(	98133	 ),
(	98158	 ),
(	98182	 ),
(	98206	 ),
(	98230	 ),
(	98255	 ),
(	98279	 ),
(	98303	 ),
(	98327	 ),
(	98352	 ),
(	98376	 ),
(	98400	 ),
(	98424	 ),
(	98448	 ),
(	98473	 ),
(	98497	 ),
(	98521	 ),
(	98545	 ),
(	98570	 ),
(	98594	 ),
(	98618	 ),
(	98642	 ),
(	98667	 ),
(	98691	 ),
(	98715	 ),
(	98739	 ),
(	98764	 ),
(	98788	 ),
(	98812	 ),
(	98836	 ),
(	98861	 ),
(	98885	 ),
(	98909	 ),
(	98933	 ),
(	98958	 ),
(	98982	 ),
(	99006	 ),
(	99030	 ),
(	99055	 ),
(	99079	 ),
(	99103	 ),
(	99127	 ),
(	99152	 ),
(	99176	 ),
(	99200	 ),
(	99224	 ),
(	99248	 ),
(	99273	 ),
(	99297	 ),
(	99321	 ),
(	99345	 ),
(	99370	 ),
(	99394	 ),
(	99418	 ),
(	99442	 ),
(	99467	 ),
(	99491	 ),
(	99515	 ),
(	99539	 ),
(	99564	 ),
(	99588	 ),
(	99612	 ),
(	99636	 ),
(	99661	 ),
(	99685	 ),
(	99709	 ),
(	99733	 ),
(	99758	 ),
(	99782	 ),
(	99806	 ),
(	99830	 ),
(	99855	 ),
(	99879	 ),
(	99903	 ),
(	99927	 ),
(	99952	 ),
(	99976	 ),
(	100000	 )
);





begin
	
	determine_limit: process (clk, distance) is
	begin
		if rising_edge(clk) then
			if to_integer(unsigned(distance)) > 3300 then
				counter_limit <= to_unsigned(100000, counter_limit'length);
			elsif to_integer(unsigned(distance)) < 0 then
				counter_limit <= to_unsigned(20000, counter_limit'length);
			else
				counter_limit <= to_unsigned(d2count(to_integer(unsigned(distance))),counter_limit'length);
			end if;
		end if;		
	end process;
	
	
	count: process (clk, reset) is
	begin		
		if rising_edge(clk) then
			if reset = '1' then
				counter <= to_unsigned(0, counter_limit'length);
			end if;
		
			counter <= counter + 1;
			
			if (counter > counter_limit) then
				counter <= to_unsigned(0, counter_limit'length);
			end if;
		end if;
	end process;
	

	produce_pwm : process(counter_limit, counter, reset)
   begin
		if reset = '1' then
			dac_out <= '0';
		else
			if (counter < (counter_limit / 2)) then  -- Potential issue unsigned(counter_limit)?
			  dac_out <= '0';
			else 
			  dac_out <= '1';
			end if;
		end if;
	end process;
				
end behavior;
